module our(clk,reset,read_base,write_base,num_read,read_size_input,read_ready,write_ready,read_data,
			read_enable,write_enable,finish_read,finish_write,read_addr,write_addr,write_size,read_size_output,write_data,done);
    input wire clk;
    input wire reset;
    input wire[63:0] read_base;
	input wire[63:0] write_base;
	input wire[63:0] num_read;
	input wire[63:0] read_size_input;
	input wire[63:0] read_ready;
	input wire[63:0] write_ready;
	input wire[63:0] read_data;
    output wire read_enable;
	output wire write_enable;
	output wire finish_read;
	output wire finish_write;
    output wire done;
	output wire[63:0] read_addr;
	output wire[63:0] write_addr;
	output wire[63:0] write_size;
	output wire[63:0] read_size_output;
    output wire[63:0] write_data;

	reg[63:0] read_cnt;
	reg[63:0] write_cnt;
	reg[63:0] state;
    reg r_read_enable;
	reg r_write_enable;
	reg r_finish_read;
	reg r_finish_write;
    reg r_done;
	reg[63:0] r_read_addr;
	reg[63:0] r_write_addr;
	reg[63:0] r_write_size;
	reg[63:0] r_read_size_output;
    //reg[63:0] r_read_data;
    reg[63:0] r_write_data;
	reg[63:0] tmp[0:201];
	reg[63:0] ans[0:201];
    assign read_enable=r_read_enable;
	assign write_enable=r_write_enable;
	assign finish_read=r_finish_read;
	assign finish_write=r_finish_write;
	assign read_addr=r_read_addr;
	assign write_addr=r_write_addr;
	assign write_size=r_write_size;
	assign read_size_output=r_read_size_output;
    assign write_data=r_write_data;
    assign done=r_done;




	parameter IDLE = 64'd0;
	parameter READY_READ = 64'd1;
	parameter WAIT_READ = 64'd2;
	parameter DEAL_READ = 64'd3;
	parameter FINISH = 64'd4;
	parameter READY_WRITE = 64'd5;
	parameter WAIT_WRITE = 64'd6;
    parameter DEAL_WRITE = 64'd7;
	parameter SUSPEND = 64'd8;
    parameter LOOP = 64'd9;
    parameter HANDLING = 64'd10;

    always @(posedge reset or posedge clk)
    begin
        if (reset)
        begin
            state<=IDLE;
            read_cnt<=0;
            write_cnt<=0;
            r_read_enable<=0;
            r_write_enable<=0;
            r_finish_read<=0;
            r_finish_write<=0;
            r_read_addr<=0;
            r_write_addr<=0;
            r_write_size<=0;
            r_read_size_output<=0;
            r_done<=0;
        end
        else
        begin
            if (state == IDLE)
            begin
                state<=WAIT_READ;
                r_read_addr<=read_base;
                r_read_size_output<=read_size_input;
                r_read_enable<=1;
            end
            else if (state == WAIT_READ)
            begin
                r_finish_read<=0;
                if (read_ready == 1)
                begin
                    tmp[read_cnt[7:0]]<=read_data;
                    state<= DEAL_READ;
                end
            end
            else if (state == DEAL_READ)
            begin
                if (read_cnt + 1 < num_read)
                begin
                    read_cnt<=read_cnt+1;
                    r_read_addr<=r_read_addr+read_size_input;
                    state<=WAIT_READ;
                    r_finish_read<=1;
                end
                else
                begin
                    state<=HANDLING;
                    r_read_enable<=0;
                    r_finish_read<=0;
                end
            end
            else if (state == HANDLING)
            begin
				ans[0]<=tmp[0]*tmp[100];
				ans[1]<=tmp[0]*tmp[101]+tmp[1]*tmp[100];
				ans[2]<=tmp[0]*tmp[102]+tmp[1]*tmp[101]+tmp[2]*tmp[100];
				ans[3]<=tmp[0]*tmp[103]+tmp[1]*tmp[102]+tmp[2]*tmp[101]+tmp[3]*tmp[100];
				ans[4]<=tmp[0]*tmp[104]+tmp[1]*tmp[103]+tmp[2]*tmp[102]+tmp[3]*tmp[101]+tmp[4]*tmp[100];
				ans[5]<=tmp[0]*tmp[105]+tmp[1]*tmp[104]+tmp[2]*tmp[103]+tmp[3]*tmp[102]+tmp[4]*tmp[101]+tmp[5]*tmp[100];
				ans[6]<=tmp[0]*tmp[106]+tmp[1]*tmp[105]+tmp[2]*tmp[104]+tmp[3]*tmp[103]+tmp[4]*tmp[102]+tmp[5]*tmp[101]+tmp[6]*tmp[100];
				ans[7]<=tmp[0]*tmp[107]+tmp[1]*tmp[106]+tmp[2]*tmp[105]+tmp[3]*tmp[104]+tmp[4]*tmp[103]+tmp[5]*tmp[102]+tmp[6]*tmp[101]+tmp[7]*tmp[100];
				ans[8]<=tmp[0]*tmp[108]+tmp[1]*tmp[107]+tmp[2]*tmp[106]+tmp[3]*tmp[105]+tmp[4]*tmp[104]+tmp[5]*tmp[103]+tmp[6]*tmp[102]+tmp[7]*tmp[101]+tmp[8]*tmp[100];
				ans[9]<=tmp[0]*tmp[109]+tmp[1]*tmp[108]+tmp[2]*tmp[107]+tmp[3]*tmp[106]+tmp[4]*tmp[105]+tmp[5]*tmp[104]+tmp[6]*tmp[103]+tmp[7]*tmp[102]+tmp[8]*tmp[101]+tmp[9]*tmp[100];
				ans[10]<=tmp[0]*tmp[110]+tmp[1]*tmp[109]+tmp[2]*tmp[108]+tmp[3]*tmp[107]+tmp[4]*tmp[106]+tmp[5]*tmp[105]+tmp[6]*tmp[104]+tmp[7]*tmp[103]+tmp[8]*tmp[102]+tmp[9]*tmp[101]+tmp[10]*tmp[100];
				ans[11]<=tmp[0]*tmp[111]+tmp[1]*tmp[110]+tmp[2]*tmp[109]+tmp[3]*tmp[108]+tmp[4]*tmp[107]+tmp[5]*tmp[106]+tmp[6]*tmp[105]+tmp[7]*tmp[104]+tmp[8]*tmp[103]+tmp[9]*tmp[102]+tmp[10]*tmp[101]+tmp[11]*tmp[100];
				ans[12]<=tmp[0]*tmp[112]+tmp[1]*tmp[111]+tmp[2]*tmp[110]+tmp[3]*tmp[109]+tmp[4]*tmp[108]+tmp[5]*tmp[107]+tmp[6]*tmp[106]+tmp[7]*tmp[105]+tmp[8]*tmp[104]+tmp[9]*tmp[103]+tmp[10]*tmp[102]+tmp[11]*tmp[101]+tmp[12]*tmp[100];
				ans[13]<=tmp[0]*tmp[113]+tmp[1]*tmp[112]+tmp[2]*tmp[111]+tmp[3]*tmp[110]+tmp[4]*tmp[109]+tmp[5]*tmp[108]+tmp[6]*tmp[107]+tmp[7]*tmp[106]+tmp[8]*tmp[105]+tmp[9]*tmp[104]+tmp[10]*tmp[103]+tmp[11]*tmp[102]+tmp[12]*tmp[101]+tmp[13]*tmp[100];
				ans[14]<=tmp[0]*tmp[114]+tmp[1]*tmp[113]+tmp[2]*tmp[112]+tmp[3]*tmp[111]+tmp[4]*tmp[110]+tmp[5]*tmp[109]+tmp[6]*tmp[108]+tmp[7]*tmp[107]+tmp[8]*tmp[106]+tmp[9]*tmp[105]+tmp[10]*tmp[104]+tmp[11]*tmp[103]+tmp[12]*tmp[102]+tmp[13]*tmp[101]+tmp[14]*tmp[100];
				ans[15]<=tmp[0]*tmp[115]+tmp[1]*tmp[114]+tmp[2]*tmp[113]+tmp[3]*tmp[112]+tmp[4]*tmp[111]+tmp[5]*tmp[110]+tmp[6]*tmp[109]+tmp[7]*tmp[108]+tmp[8]*tmp[107]+tmp[9]*tmp[106]+tmp[10]*tmp[105]+tmp[11]*tmp[104]+tmp[12]*tmp[103]+tmp[13]*tmp[102]+tmp[14]*tmp[101]+tmp[15]*tmp[100];
				ans[16]<=tmp[0]*tmp[116]+tmp[1]*tmp[115]+tmp[2]*tmp[114]+tmp[3]*tmp[113]+tmp[4]*tmp[112]+tmp[5]*tmp[111]+tmp[6]*tmp[110]+tmp[7]*tmp[109]+tmp[8]*tmp[108]+tmp[9]*tmp[107]+tmp[10]*tmp[106]+tmp[11]*tmp[105]+tmp[12]*tmp[104]+tmp[13]*tmp[103]+tmp[14]*tmp[102]+tmp[15]*tmp[101]+tmp[16]*tmp[100];
				ans[17]<=tmp[0]*tmp[117]+tmp[1]*tmp[116]+tmp[2]*tmp[115]+tmp[3]*tmp[114]+tmp[4]*tmp[113]+tmp[5]*tmp[112]+tmp[6]*tmp[111]+tmp[7]*tmp[110]+tmp[8]*tmp[109]+tmp[9]*tmp[108]+tmp[10]*tmp[107]+tmp[11]*tmp[106]+tmp[12]*tmp[105]+tmp[13]*tmp[104]+tmp[14]*tmp[103]+tmp[15]*tmp[102]+tmp[16]*tmp[101]+tmp[17]*tmp[100];
				ans[18]<=tmp[0]*tmp[118]+tmp[1]*tmp[117]+tmp[2]*tmp[116]+tmp[3]*tmp[115]+tmp[4]*tmp[114]+tmp[5]*tmp[113]+tmp[6]*tmp[112]+tmp[7]*tmp[111]+tmp[8]*tmp[110]+tmp[9]*tmp[109]+tmp[10]*tmp[108]+tmp[11]*tmp[107]+tmp[12]*tmp[106]+tmp[13]*tmp[105]+tmp[14]*tmp[104]+tmp[15]*tmp[103]+tmp[16]*tmp[102]+tmp[17]*tmp[101]+tmp[18]*tmp[100];
				ans[19]<=tmp[0]*tmp[119]+tmp[1]*tmp[118]+tmp[2]*tmp[117]+tmp[3]*tmp[116]+tmp[4]*tmp[115]+tmp[5]*tmp[114]+tmp[6]*tmp[113]+tmp[7]*tmp[112]+tmp[8]*tmp[111]+tmp[9]*tmp[110]+tmp[10]*tmp[109]+tmp[11]*tmp[108]+tmp[12]*tmp[107]+tmp[13]*tmp[106]+tmp[14]*tmp[105]+tmp[15]*tmp[104]+tmp[16]*tmp[103]+tmp[17]*tmp[102]+tmp[18]*tmp[101]+tmp[19]*tmp[100];
				ans[20]<=tmp[0]*tmp[120]+tmp[1]*tmp[119]+tmp[2]*tmp[118]+tmp[3]*tmp[117]+tmp[4]*tmp[116]+tmp[5]*tmp[115]+tmp[6]*tmp[114]+tmp[7]*tmp[113]+tmp[8]*tmp[112]+tmp[9]*tmp[111]+tmp[10]*tmp[110]+tmp[11]*tmp[109]+tmp[12]*tmp[108]+tmp[13]*tmp[107]+tmp[14]*tmp[106]+tmp[15]*tmp[105]+tmp[16]*tmp[104]+tmp[17]*tmp[103]+tmp[18]*tmp[102]+tmp[19]*tmp[101]+tmp[20]*tmp[100];
				ans[21]<=tmp[0]*tmp[121]+tmp[1]*tmp[120]+tmp[2]*tmp[119]+tmp[3]*tmp[118]+tmp[4]*tmp[117]+tmp[5]*tmp[116]+tmp[6]*tmp[115]+tmp[7]*tmp[114]+tmp[8]*tmp[113]+tmp[9]*tmp[112]+tmp[10]*tmp[111]+tmp[11]*tmp[110]+tmp[12]*tmp[109]+tmp[13]*tmp[108]+tmp[14]*tmp[107]+tmp[15]*tmp[106]+tmp[16]*tmp[105]+tmp[17]*tmp[104]+tmp[18]*tmp[103]+tmp[19]*tmp[102]+tmp[20]*tmp[101]+tmp[21]*tmp[100];
				ans[22]<=tmp[0]*tmp[122]+tmp[1]*tmp[121]+tmp[2]*tmp[120]+tmp[3]*tmp[119]+tmp[4]*tmp[118]+tmp[5]*tmp[117]+tmp[6]*tmp[116]+tmp[7]*tmp[115]+tmp[8]*tmp[114]+tmp[9]*tmp[113]+tmp[10]*tmp[112]+tmp[11]*tmp[111]+tmp[12]*tmp[110]+tmp[13]*tmp[109]+tmp[14]*tmp[108]+tmp[15]*tmp[107]+tmp[16]*tmp[106]+tmp[17]*tmp[105]+tmp[18]*tmp[104]+tmp[19]*tmp[103]+tmp[20]*tmp[102]+tmp[21]*tmp[101]+tmp[22]*tmp[100];
				ans[23]<=tmp[0]*tmp[123]+tmp[1]*tmp[122]+tmp[2]*tmp[121]+tmp[3]*tmp[120]+tmp[4]*tmp[119]+tmp[5]*tmp[118]+tmp[6]*tmp[117]+tmp[7]*tmp[116]+tmp[8]*tmp[115]+tmp[9]*tmp[114]+tmp[10]*tmp[113]+tmp[11]*tmp[112]+tmp[12]*tmp[111]+tmp[13]*tmp[110]+tmp[14]*tmp[109]+tmp[15]*tmp[108]+tmp[16]*tmp[107]+tmp[17]*tmp[106]+tmp[18]*tmp[105]+tmp[19]*tmp[104]+tmp[20]*tmp[103]+tmp[21]*tmp[102]+tmp[22]*tmp[101]+tmp[23]*tmp[100];
				ans[24]<=tmp[0]*tmp[124]+tmp[1]*tmp[123]+tmp[2]*tmp[122]+tmp[3]*tmp[121]+tmp[4]*tmp[120]+tmp[5]*tmp[119]+tmp[6]*tmp[118]+tmp[7]*tmp[117]+tmp[8]*tmp[116]+tmp[9]*tmp[115]+tmp[10]*tmp[114]+tmp[11]*tmp[113]+tmp[12]*tmp[112]+tmp[13]*tmp[111]+tmp[14]*tmp[110]+tmp[15]*tmp[109]+tmp[16]*tmp[108]+tmp[17]*tmp[107]+tmp[18]*tmp[106]+tmp[19]*tmp[105]+tmp[20]*tmp[104]+tmp[21]*tmp[103]+tmp[22]*tmp[102]+tmp[23]*tmp[101]+tmp[24]*tmp[100];
				ans[25]<=tmp[0]*tmp[125]+tmp[1]*tmp[124]+tmp[2]*tmp[123]+tmp[3]*tmp[122]+tmp[4]*tmp[121]+tmp[5]*tmp[120]+tmp[6]*tmp[119]+tmp[7]*tmp[118]+tmp[8]*tmp[117]+tmp[9]*tmp[116]+tmp[10]*tmp[115]+tmp[11]*tmp[114]+tmp[12]*tmp[113]+tmp[13]*tmp[112]+tmp[14]*tmp[111]+tmp[15]*tmp[110]+tmp[16]*tmp[109]+tmp[17]*tmp[108]+tmp[18]*tmp[107]+tmp[19]*tmp[106]+tmp[20]*tmp[105]+tmp[21]*tmp[104]+tmp[22]*tmp[103]+tmp[23]*tmp[102]+tmp[24]*tmp[101]+tmp[25]*tmp[100];
				ans[26]<=tmp[0]*tmp[126]+tmp[1]*tmp[125]+tmp[2]*tmp[124]+tmp[3]*tmp[123]+tmp[4]*tmp[122]+tmp[5]*tmp[121]+tmp[6]*tmp[120]+tmp[7]*tmp[119]+tmp[8]*tmp[118]+tmp[9]*tmp[117]+tmp[10]*tmp[116]+tmp[11]*tmp[115]+tmp[12]*tmp[114]+tmp[13]*tmp[113]+tmp[14]*tmp[112]+tmp[15]*tmp[111]+tmp[16]*tmp[110]+tmp[17]*tmp[109]+tmp[18]*tmp[108]+tmp[19]*tmp[107]+tmp[20]*tmp[106]+tmp[21]*tmp[105]+tmp[22]*tmp[104]+tmp[23]*tmp[103]+tmp[24]*tmp[102]+tmp[25]*tmp[101]+tmp[26]*tmp[100];
				ans[27]<=tmp[0]*tmp[127]+tmp[1]*tmp[126]+tmp[2]*tmp[125]+tmp[3]*tmp[124]+tmp[4]*tmp[123]+tmp[5]*tmp[122]+tmp[6]*tmp[121]+tmp[7]*tmp[120]+tmp[8]*tmp[119]+tmp[9]*tmp[118]+tmp[10]*tmp[117]+tmp[11]*tmp[116]+tmp[12]*tmp[115]+tmp[13]*tmp[114]+tmp[14]*tmp[113]+tmp[15]*tmp[112]+tmp[16]*tmp[111]+tmp[17]*tmp[110]+tmp[18]*tmp[109]+tmp[19]*tmp[108]+tmp[20]*tmp[107]+tmp[21]*tmp[106]+tmp[22]*tmp[105]+tmp[23]*tmp[104]+tmp[24]*tmp[103]+tmp[25]*tmp[102]+tmp[26]*tmp[101]+tmp[27]*tmp[100];
				ans[28]<=tmp[0]*tmp[128]+tmp[1]*tmp[127]+tmp[2]*tmp[126]+tmp[3]*tmp[125]+tmp[4]*tmp[124]+tmp[5]*tmp[123]+tmp[6]*tmp[122]+tmp[7]*tmp[121]+tmp[8]*tmp[120]+tmp[9]*tmp[119]+tmp[10]*tmp[118]+tmp[11]*tmp[117]+tmp[12]*tmp[116]+tmp[13]*tmp[115]+tmp[14]*tmp[114]+tmp[15]*tmp[113]+tmp[16]*tmp[112]+tmp[17]*tmp[111]+tmp[18]*tmp[110]+tmp[19]*tmp[109]+tmp[20]*tmp[108]+tmp[21]*tmp[107]+tmp[22]*tmp[106]+tmp[23]*tmp[105]+tmp[24]*tmp[104]+tmp[25]*tmp[103]+tmp[26]*tmp[102]+tmp[27]*tmp[101]+tmp[28]*tmp[100];
				ans[29]<=tmp[0]*tmp[129]+tmp[1]*tmp[128]+tmp[2]*tmp[127]+tmp[3]*tmp[126]+tmp[4]*tmp[125]+tmp[5]*tmp[124]+tmp[6]*tmp[123]+tmp[7]*tmp[122]+tmp[8]*tmp[121]+tmp[9]*tmp[120]+tmp[10]*tmp[119]+tmp[11]*tmp[118]+tmp[12]*tmp[117]+tmp[13]*tmp[116]+tmp[14]*tmp[115]+tmp[15]*tmp[114]+tmp[16]*tmp[113]+tmp[17]*tmp[112]+tmp[18]*tmp[111]+tmp[19]*tmp[110]+tmp[20]*tmp[109]+tmp[21]*tmp[108]+tmp[22]*tmp[107]+tmp[23]*tmp[106]+tmp[24]*tmp[105]+tmp[25]*tmp[104]+tmp[26]*tmp[103]+tmp[27]*tmp[102]+tmp[28]*tmp[101]+tmp[29]*tmp[100];
				ans[30]<=tmp[0]*tmp[130]+tmp[1]*tmp[129]+tmp[2]*tmp[128]+tmp[3]*tmp[127]+tmp[4]*tmp[126]+tmp[5]*tmp[125]+tmp[6]*tmp[124]+tmp[7]*tmp[123]+tmp[8]*tmp[122]+tmp[9]*tmp[121]+tmp[10]*tmp[120]+tmp[11]*tmp[119]+tmp[12]*tmp[118]+tmp[13]*tmp[117]+tmp[14]*tmp[116]+tmp[15]*tmp[115]+tmp[16]*tmp[114]+tmp[17]*tmp[113]+tmp[18]*tmp[112]+tmp[19]*tmp[111]+tmp[20]*tmp[110]+tmp[21]*tmp[109]+tmp[22]*tmp[108]+tmp[23]*tmp[107]+tmp[24]*tmp[106]+tmp[25]*tmp[105]+tmp[26]*tmp[104]+tmp[27]*tmp[103]+tmp[28]*tmp[102]+tmp[29]*tmp[101]+tmp[30]*tmp[100];
				ans[31]<=tmp[0]*tmp[131]+tmp[1]*tmp[130]+tmp[2]*tmp[129]+tmp[3]*tmp[128]+tmp[4]*tmp[127]+tmp[5]*tmp[126]+tmp[6]*tmp[125]+tmp[7]*tmp[124]+tmp[8]*tmp[123]+tmp[9]*tmp[122]+tmp[10]*tmp[121]+tmp[11]*tmp[120]+tmp[12]*tmp[119]+tmp[13]*tmp[118]+tmp[14]*tmp[117]+tmp[15]*tmp[116]+tmp[16]*tmp[115]+tmp[17]*tmp[114]+tmp[18]*tmp[113]+tmp[19]*tmp[112]+tmp[20]*tmp[111]+tmp[21]*tmp[110]+tmp[22]*tmp[109]+tmp[23]*tmp[108]+tmp[24]*tmp[107]+tmp[25]*tmp[106]+tmp[26]*tmp[105]+tmp[27]*tmp[104]+tmp[28]*tmp[103]+tmp[29]*tmp[102]+tmp[30]*tmp[101]+tmp[31]*tmp[100];
				ans[32]<=tmp[0]*tmp[132]+tmp[1]*tmp[131]+tmp[2]*tmp[130]+tmp[3]*tmp[129]+tmp[4]*tmp[128]+tmp[5]*tmp[127]+tmp[6]*tmp[126]+tmp[7]*tmp[125]+tmp[8]*tmp[124]+tmp[9]*tmp[123]+tmp[10]*tmp[122]+tmp[11]*tmp[121]+tmp[12]*tmp[120]+tmp[13]*tmp[119]+tmp[14]*tmp[118]+tmp[15]*tmp[117]+tmp[16]*tmp[116]+tmp[17]*tmp[115]+tmp[18]*tmp[114]+tmp[19]*tmp[113]+tmp[20]*tmp[112]+tmp[21]*tmp[111]+tmp[22]*tmp[110]+tmp[23]*tmp[109]+tmp[24]*tmp[108]+tmp[25]*tmp[107]+tmp[26]*tmp[106]+tmp[27]*tmp[105]+tmp[28]*tmp[104]+tmp[29]*tmp[103]+tmp[30]*tmp[102]+tmp[31]*tmp[101]+tmp[32]*tmp[100];
				ans[33]<=tmp[0]*tmp[133]+tmp[1]*tmp[132]+tmp[2]*tmp[131]+tmp[3]*tmp[130]+tmp[4]*tmp[129]+tmp[5]*tmp[128]+tmp[6]*tmp[127]+tmp[7]*tmp[126]+tmp[8]*tmp[125]+tmp[9]*tmp[124]+tmp[10]*tmp[123]+tmp[11]*tmp[122]+tmp[12]*tmp[121]+tmp[13]*tmp[120]+tmp[14]*tmp[119]+tmp[15]*tmp[118]+tmp[16]*tmp[117]+tmp[17]*tmp[116]+tmp[18]*tmp[115]+tmp[19]*tmp[114]+tmp[20]*tmp[113]+tmp[21]*tmp[112]+tmp[22]*tmp[111]+tmp[23]*tmp[110]+tmp[24]*tmp[109]+tmp[25]*tmp[108]+tmp[26]*tmp[107]+tmp[27]*tmp[106]+tmp[28]*tmp[105]+tmp[29]*tmp[104]+tmp[30]*tmp[103]+tmp[31]*tmp[102]+tmp[32]*tmp[101]+tmp[33]*tmp[100];
				ans[34]<=tmp[0]*tmp[134]+tmp[1]*tmp[133]+tmp[2]*tmp[132]+tmp[3]*tmp[131]+tmp[4]*tmp[130]+tmp[5]*tmp[129]+tmp[6]*tmp[128]+tmp[7]*tmp[127]+tmp[8]*tmp[126]+tmp[9]*tmp[125]+tmp[10]*tmp[124]+tmp[11]*tmp[123]+tmp[12]*tmp[122]+tmp[13]*tmp[121]+tmp[14]*tmp[120]+tmp[15]*tmp[119]+tmp[16]*tmp[118]+tmp[17]*tmp[117]+tmp[18]*tmp[116]+tmp[19]*tmp[115]+tmp[20]*tmp[114]+tmp[21]*tmp[113]+tmp[22]*tmp[112]+tmp[23]*tmp[111]+tmp[24]*tmp[110]+tmp[25]*tmp[109]+tmp[26]*tmp[108]+tmp[27]*tmp[107]+tmp[28]*tmp[106]+tmp[29]*tmp[105]+tmp[30]*tmp[104]+tmp[31]*tmp[103]+tmp[32]*tmp[102]+tmp[33]*tmp[101]+tmp[34]*tmp[100];
				ans[35]<=tmp[0]*tmp[135]+tmp[1]*tmp[134]+tmp[2]*tmp[133]+tmp[3]*tmp[132]+tmp[4]*tmp[131]+tmp[5]*tmp[130]+tmp[6]*tmp[129]+tmp[7]*tmp[128]+tmp[8]*tmp[127]+tmp[9]*tmp[126]+tmp[10]*tmp[125]+tmp[11]*tmp[124]+tmp[12]*tmp[123]+tmp[13]*tmp[122]+tmp[14]*tmp[121]+tmp[15]*tmp[120]+tmp[16]*tmp[119]+tmp[17]*tmp[118]+tmp[18]*tmp[117]+tmp[19]*tmp[116]+tmp[20]*tmp[115]+tmp[21]*tmp[114]+tmp[22]*tmp[113]+tmp[23]*tmp[112]+tmp[24]*tmp[111]+tmp[25]*tmp[110]+tmp[26]*tmp[109]+tmp[27]*tmp[108]+tmp[28]*tmp[107]+tmp[29]*tmp[106]+tmp[30]*tmp[105]+tmp[31]*tmp[104]+tmp[32]*tmp[103]+tmp[33]*tmp[102]+tmp[34]*tmp[101]+tmp[35]*tmp[100];
				ans[36]<=tmp[0]*tmp[136]+tmp[1]*tmp[135]+tmp[2]*tmp[134]+tmp[3]*tmp[133]+tmp[4]*tmp[132]+tmp[5]*tmp[131]+tmp[6]*tmp[130]+tmp[7]*tmp[129]+tmp[8]*tmp[128]+tmp[9]*tmp[127]+tmp[10]*tmp[126]+tmp[11]*tmp[125]+tmp[12]*tmp[124]+tmp[13]*tmp[123]+tmp[14]*tmp[122]+tmp[15]*tmp[121]+tmp[16]*tmp[120]+tmp[17]*tmp[119]+tmp[18]*tmp[118]+tmp[19]*tmp[117]+tmp[20]*tmp[116]+tmp[21]*tmp[115]+tmp[22]*tmp[114]+tmp[23]*tmp[113]+tmp[24]*tmp[112]+tmp[25]*tmp[111]+tmp[26]*tmp[110]+tmp[27]*tmp[109]+tmp[28]*tmp[108]+tmp[29]*tmp[107]+tmp[30]*tmp[106]+tmp[31]*tmp[105]+tmp[32]*tmp[104]+tmp[33]*tmp[103]+tmp[34]*tmp[102]+tmp[35]*tmp[101]+tmp[36]*tmp[100];
				ans[37]<=tmp[0]*tmp[137]+tmp[1]*tmp[136]+tmp[2]*tmp[135]+tmp[3]*tmp[134]+tmp[4]*tmp[133]+tmp[5]*tmp[132]+tmp[6]*tmp[131]+tmp[7]*tmp[130]+tmp[8]*tmp[129]+tmp[9]*tmp[128]+tmp[10]*tmp[127]+tmp[11]*tmp[126]+tmp[12]*tmp[125]+tmp[13]*tmp[124]+tmp[14]*tmp[123]+tmp[15]*tmp[122]+tmp[16]*tmp[121]+tmp[17]*tmp[120]+tmp[18]*tmp[119]+tmp[19]*tmp[118]+tmp[20]*tmp[117]+tmp[21]*tmp[116]+tmp[22]*tmp[115]+tmp[23]*tmp[114]+tmp[24]*tmp[113]+tmp[25]*tmp[112]+tmp[26]*tmp[111]+tmp[27]*tmp[110]+tmp[28]*tmp[109]+tmp[29]*tmp[108]+tmp[30]*tmp[107]+tmp[31]*tmp[106]+tmp[32]*tmp[105]+tmp[33]*tmp[104]+tmp[34]*tmp[103]+tmp[35]*tmp[102]+tmp[36]*tmp[101]+tmp[37]*tmp[100];
				ans[38]<=tmp[0]*tmp[138]+tmp[1]*tmp[137]+tmp[2]*tmp[136]+tmp[3]*tmp[135]+tmp[4]*tmp[134]+tmp[5]*tmp[133]+tmp[6]*tmp[132]+tmp[7]*tmp[131]+tmp[8]*tmp[130]+tmp[9]*tmp[129]+tmp[10]*tmp[128]+tmp[11]*tmp[127]+tmp[12]*tmp[126]+tmp[13]*tmp[125]+tmp[14]*tmp[124]+tmp[15]*tmp[123]+tmp[16]*tmp[122]+tmp[17]*tmp[121]+tmp[18]*tmp[120]+tmp[19]*tmp[119]+tmp[20]*tmp[118]+tmp[21]*tmp[117]+tmp[22]*tmp[116]+tmp[23]*tmp[115]+tmp[24]*tmp[114]+tmp[25]*tmp[113]+tmp[26]*tmp[112]+tmp[27]*tmp[111]+tmp[28]*tmp[110]+tmp[29]*tmp[109]+tmp[30]*tmp[108]+tmp[31]*tmp[107]+tmp[32]*tmp[106]+tmp[33]*tmp[105]+tmp[34]*tmp[104]+tmp[35]*tmp[103]+tmp[36]*tmp[102]+tmp[37]*tmp[101]+tmp[38]*tmp[100];
				ans[39]<=tmp[0]*tmp[139]+tmp[1]*tmp[138]+tmp[2]*tmp[137]+tmp[3]*tmp[136]+tmp[4]*tmp[135]+tmp[5]*tmp[134]+tmp[6]*tmp[133]+tmp[7]*tmp[132]+tmp[8]*tmp[131]+tmp[9]*tmp[130]+tmp[10]*tmp[129]+tmp[11]*tmp[128]+tmp[12]*tmp[127]+tmp[13]*tmp[126]+tmp[14]*tmp[125]+tmp[15]*tmp[124]+tmp[16]*tmp[123]+tmp[17]*tmp[122]+tmp[18]*tmp[121]+tmp[19]*tmp[120]+tmp[20]*tmp[119]+tmp[21]*tmp[118]+tmp[22]*tmp[117]+tmp[23]*tmp[116]+tmp[24]*tmp[115]+tmp[25]*tmp[114]+tmp[26]*tmp[113]+tmp[27]*tmp[112]+tmp[28]*tmp[111]+tmp[29]*tmp[110]+tmp[30]*tmp[109]+tmp[31]*tmp[108]+tmp[32]*tmp[107]+tmp[33]*tmp[106]+tmp[34]*tmp[105]+tmp[35]*tmp[104]+tmp[36]*tmp[103]+tmp[37]*tmp[102]+tmp[38]*tmp[101]+tmp[39]*tmp[100];
				ans[40]<=tmp[0]*tmp[140]+tmp[1]*tmp[139]+tmp[2]*tmp[138]+tmp[3]*tmp[137]+tmp[4]*tmp[136]+tmp[5]*tmp[135]+tmp[6]*tmp[134]+tmp[7]*tmp[133]+tmp[8]*tmp[132]+tmp[9]*tmp[131]+tmp[10]*tmp[130]+tmp[11]*tmp[129]+tmp[12]*tmp[128]+tmp[13]*tmp[127]+tmp[14]*tmp[126]+tmp[15]*tmp[125]+tmp[16]*tmp[124]+tmp[17]*tmp[123]+tmp[18]*tmp[122]+tmp[19]*tmp[121]+tmp[20]*tmp[120]+tmp[21]*tmp[119]+tmp[22]*tmp[118]+tmp[23]*tmp[117]+tmp[24]*tmp[116]+tmp[25]*tmp[115]+tmp[26]*tmp[114]+tmp[27]*tmp[113]+tmp[28]*tmp[112]+tmp[29]*tmp[111]+tmp[30]*tmp[110]+tmp[31]*tmp[109]+tmp[32]*tmp[108]+tmp[33]*tmp[107]+tmp[34]*tmp[106]+tmp[35]*tmp[105]+tmp[36]*tmp[104]+tmp[37]*tmp[103]+tmp[38]*tmp[102]+tmp[39]*tmp[101]+tmp[40]*tmp[100];
				ans[41]<=tmp[0]*tmp[141]+tmp[1]*tmp[140]+tmp[2]*tmp[139]+tmp[3]*tmp[138]+tmp[4]*tmp[137]+tmp[5]*tmp[136]+tmp[6]*tmp[135]+tmp[7]*tmp[134]+tmp[8]*tmp[133]+tmp[9]*tmp[132]+tmp[10]*tmp[131]+tmp[11]*tmp[130]+tmp[12]*tmp[129]+tmp[13]*tmp[128]+tmp[14]*tmp[127]+tmp[15]*tmp[126]+tmp[16]*tmp[125]+tmp[17]*tmp[124]+tmp[18]*tmp[123]+tmp[19]*tmp[122]+tmp[20]*tmp[121]+tmp[21]*tmp[120]+tmp[22]*tmp[119]+tmp[23]*tmp[118]+tmp[24]*tmp[117]+tmp[25]*tmp[116]+tmp[26]*tmp[115]+tmp[27]*tmp[114]+tmp[28]*tmp[113]+tmp[29]*tmp[112]+tmp[30]*tmp[111]+tmp[31]*tmp[110]+tmp[32]*tmp[109]+tmp[33]*tmp[108]+tmp[34]*tmp[107]+tmp[35]*tmp[106]+tmp[36]*tmp[105]+tmp[37]*tmp[104]+tmp[38]*tmp[103]+tmp[39]*tmp[102]+tmp[40]*tmp[101]+tmp[41]*tmp[100];
				ans[42]<=tmp[0]*tmp[142]+tmp[1]*tmp[141]+tmp[2]*tmp[140]+tmp[3]*tmp[139]+tmp[4]*tmp[138]+tmp[5]*tmp[137]+tmp[6]*tmp[136]+tmp[7]*tmp[135]+tmp[8]*tmp[134]+tmp[9]*tmp[133]+tmp[10]*tmp[132]+tmp[11]*tmp[131]+tmp[12]*tmp[130]+tmp[13]*tmp[129]+tmp[14]*tmp[128]+tmp[15]*tmp[127]+tmp[16]*tmp[126]+tmp[17]*tmp[125]+tmp[18]*tmp[124]+tmp[19]*tmp[123]+tmp[20]*tmp[122]+tmp[21]*tmp[121]+tmp[22]*tmp[120]+tmp[23]*tmp[119]+tmp[24]*tmp[118]+tmp[25]*tmp[117]+tmp[26]*tmp[116]+tmp[27]*tmp[115]+tmp[28]*tmp[114]+tmp[29]*tmp[113]+tmp[30]*tmp[112]+tmp[31]*tmp[111]+tmp[32]*tmp[110]+tmp[33]*tmp[109]+tmp[34]*tmp[108]+tmp[35]*tmp[107]+tmp[36]*tmp[106]+tmp[37]*tmp[105]+tmp[38]*tmp[104]+tmp[39]*tmp[103]+tmp[40]*tmp[102]+tmp[41]*tmp[101]+tmp[42]*tmp[100];
				ans[43]<=tmp[0]*tmp[143]+tmp[1]*tmp[142]+tmp[2]*tmp[141]+tmp[3]*tmp[140]+tmp[4]*tmp[139]+tmp[5]*tmp[138]+tmp[6]*tmp[137]+tmp[7]*tmp[136]+tmp[8]*tmp[135]+tmp[9]*tmp[134]+tmp[10]*tmp[133]+tmp[11]*tmp[132]+tmp[12]*tmp[131]+tmp[13]*tmp[130]+tmp[14]*tmp[129]+tmp[15]*tmp[128]+tmp[16]*tmp[127]+tmp[17]*tmp[126]+tmp[18]*tmp[125]+tmp[19]*tmp[124]+tmp[20]*tmp[123]+tmp[21]*tmp[122]+tmp[22]*tmp[121]+tmp[23]*tmp[120]+tmp[24]*tmp[119]+tmp[25]*tmp[118]+tmp[26]*tmp[117]+tmp[27]*tmp[116]+tmp[28]*tmp[115]+tmp[29]*tmp[114]+tmp[30]*tmp[113]+tmp[31]*tmp[112]+tmp[32]*tmp[111]+tmp[33]*tmp[110]+tmp[34]*tmp[109]+tmp[35]*tmp[108]+tmp[36]*tmp[107]+tmp[37]*tmp[106]+tmp[38]*tmp[105]+tmp[39]*tmp[104]+tmp[40]*tmp[103]+tmp[41]*tmp[102]+tmp[42]*tmp[101]+tmp[43]*tmp[100];
				ans[44]<=tmp[0]*tmp[144]+tmp[1]*tmp[143]+tmp[2]*tmp[142]+tmp[3]*tmp[141]+tmp[4]*tmp[140]+tmp[5]*tmp[139]+tmp[6]*tmp[138]+tmp[7]*tmp[137]+tmp[8]*tmp[136]+tmp[9]*tmp[135]+tmp[10]*tmp[134]+tmp[11]*tmp[133]+tmp[12]*tmp[132]+tmp[13]*tmp[131]+tmp[14]*tmp[130]+tmp[15]*tmp[129]+tmp[16]*tmp[128]+tmp[17]*tmp[127]+tmp[18]*tmp[126]+tmp[19]*tmp[125]+tmp[20]*tmp[124]+tmp[21]*tmp[123]+tmp[22]*tmp[122]+tmp[23]*tmp[121]+tmp[24]*tmp[120]+tmp[25]*tmp[119]+tmp[26]*tmp[118]+tmp[27]*tmp[117]+tmp[28]*tmp[116]+tmp[29]*tmp[115]+tmp[30]*tmp[114]+tmp[31]*tmp[113]+tmp[32]*tmp[112]+tmp[33]*tmp[111]+tmp[34]*tmp[110]+tmp[35]*tmp[109]+tmp[36]*tmp[108]+tmp[37]*tmp[107]+tmp[38]*tmp[106]+tmp[39]*tmp[105]+tmp[40]*tmp[104]+tmp[41]*tmp[103]+tmp[42]*tmp[102]+tmp[43]*tmp[101]+tmp[44]*tmp[100];
				ans[45]<=tmp[0]*tmp[145]+tmp[1]*tmp[144]+tmp[2]*tmp[143]+tmp[3]*tmp[142]+tmp[4]*tmp[141]+tmp[5]*tmp[140]+tmp[6]*tmp[139]+tmp[7]*tmp[138]+tmp[8]*tmp[137]+tmp[9]*tmp[136]+tmp[10]*tmp[135]+tmp[11]*tmp[134]+tmp[12]*tmp[133]+tmp[13]*tmp[132]+tmp[14]*tmp[131]+tmp[15]*tmp[130]+tmp[16]*tmp[129]+tmp[17]*tmp[128]+tmp[18]*tmp[127]+tmp[19]*tmp[126]+tmp[20]*tmp[125]+tmp[21]*tmp[124]+tmp[22]*tmp[123]+tmp[23]*tmp[122]+tmp[24]*tmp[121]+tmp[25]*tmp[120]+tmp[26]*tmp[119]+tmp[27]*tmp[118]+tmp[28]*tmp[117]+tmp[29]*tmp[116]+tmp[30]*tmp[115]+tmp[31]*tmp[114]+tmp[32]*tmp[113]+tmp[33]*tmp[112]+tmp[34]*tmp[111]+tmp[35]*tmp[110]+tmp[36]*tmp[109]+tmp[37]*tmp[108]+tmp[38]*tmp[107]+tmp[39]*tmp[106]+tmp[40]*tmp[105]+tmp[41]*tmp[104]+tmp[42]*tmp[103]+tmp[43]*tmp[102]+tmp[44]*tmp[101]+tmp[45]*tmp[100];
				ans[46]<=tmp[0]*tmp[146]+tmp[1]*tmp[145]+tmp[2]*tmp[144]+tmp[3]*tmp[143]+tmp[4]*tmp[142]+tmp[5]*tmp[141]+tmp[6]*tmp[140]+tmp[7]*tmp[139]+tmp[8]*tmp[138]+tmp[9]*tmp[137]+tmp[10]*tmp[136]+tmp[11]*tmp[135]+tmp[12]*tmp[134]+tmp[13]*tmp[133]+tmp[14]*tmp[132]+tmp[15]*tmp[131]+tmp[16]*tmp[130]+tmp[17]*tmp[129]+tmp[18]*tmp[128]+tmp[19]*tmp[127]+tmp[20]*tmp[126]+tmp[21]*tmp[125]+tmp[22]*tmp[124]+tmp[23]*tmp[123]+tmp[24]*tmp[122]+tmp[25]*tmp[121]+tmp[26]*tmp[120]+tmp[27]*tmp[119]+tmp[28]*tmp[118]+tmp[29]*tmp[117]+tmp[30]*tmp[116]+tmp[31]*tmp[115]+tmp[32]*tmp[114]+tmp[33]*tmp[113]+tmp[34]*tmp[112]+tmp[35]*tmp[111]+tmp[36]*tmp[110]+tmp[37]*tmp[109]+tmp[38]*tmp[108]+tmp[39]*tmp[107]+tmp[40]*tmp[106]+tmp[41]*tmp[105]+tmp[42]*tmp[104]+tmp[43]*tmp[103]+tmp[44]*tmp[102]+tmp[45]*tmp[101]+tmp[46]*tmp[100];
				ans[47]<=tmp[0]*tmp[147]+tmp[1]*tmp[146]+tmp[2]*tmp[145]+tmp[3]*tmp[144]+tmp[4]*tmp[143]+tmp[5]*tmp[142]+tmp[6]*tmp[141]+tmp[7]*tmp[140]+tmp[8]*tmp[139]+tmp[9]*tmp[138]+tmp[10]*tmp[137]+tmp[11]*tmp[136]+tmp[12]*tmp[135]+tmp[13]*tmp[134]+tmp[14]*tmp[133]+tmp[15]*tmp[132]+tmp[16]*tmp[131]+tmp[17]*tmp[130]+tmp[18]*tmp[129]+tmp[19]*tmp[128]+tmp[20]*tmp[127]+tmp[21]*tmp[126]+tmp[22]*tmp[125]+tmp[23]*tmp[124]+tmp[24]*tmp[123]+tmp[25]*tmp[122]+tmp[26]*tmp[121]+tmp[27]*tmp[120]+tmp[28]*tmp[119]+tmp[29]*tmp[118]+tmp[30]*tmp[117]+tmp[31]*tmp[116]+tmp[32]*tmp[115]+tmp[33]*tmp[114]+tmp[34]*tmp[113]+tmp[35]*tmp[112]+tmp[36]*tmp[111]+tmp[37]*tmp[110]+tmp[38]*tmp[109]+tmp[39]*tmp[108]+tmp[40]*tmp[107]+tmp[41]*tmp[106]+tmp[42]*tmp[105]+tmp[43]*tmp[104]+tmp[44]*tmp[103]+tmp[45]*tmp[102]+tmp[46]*tmp[101]+tmp[47]*tmp[100];
				ans[48]<=tmp[0]*tmp[148]+tmp[1]*tmp[147]+tmp[2]*tmp[146]+tmp[3]*tmp[145]+tmp[4]*tmp[144]+tmp[5]*tmp[143]+tmp[6]*tmp[142]+tmp[7]*tmp[141]+tmp[8]*tmp[140]+tmp[9]*tmp[139]+tmp[10]*tmp[138]+tmp[11]*tmp[137]+tmp[12]*tmp[136]+tmp[13]*tmp[135]+tmp[14]*tmp[134]+tmp[15]*tmp[133]+tmp[16]*tmp[132]+tmp[17]*tmp[131]+tmp[18]*tmp[130]+tmp[19]*tmp[129]+tmp[20]*tmp[128]+tmp[21]*tmp[127]+tmp[22]*tmp[126]+tmp[23]*tmp[125]+tmp[24]*tmp[124]+tmp[25]*tmp[123]+tmp[26]*tmp[122]+tmp[27]*tmp[121]+tmp[28]*tmp[120]+tmp[29]*tmp[119]+tmp[30]*tmp[118]+tmp[31]*tmp[117]+tmp[32]*tmp[116]+tmp[33]*tmp[115]+tmp[34]*tmp[114]+tmp[35]*tmp[113]+tmp[36]*tmp[112]+tmp[37]*tmp[111]+tmp[38]*tmp[110]+tmp[39]*tmp[109]+tmp[40]*tmp[108]+tmp[41]*tmp[107]+tmp[42]*tmp[106]+tmp[43]*tmp[105]+tmp[44]*tmp[104]+tmp[45]*tmp[103]+tmp[46]*tmp[102]+tmp[47]*tmp[101]+tmp[48]*tmp[100];
				ans[49]<=tmp[0]*tmp[149]+tmp[1]*tmp[148]+tmp[2]*tmp[147]+tmp[3]*tmp[146]+tmp[4]*tmp[145]+tmp[5]*tmp[144]+tmp[6]*tmp[143]+tmp[7]*tmp[142]+tmp[8]*tmp[141]+tmp[9]*tmp[140]+tmp[10]*tmp[139]+tmp[11]*tmp[138]+tmp[12]*tmp[137]+tmp[13]*tmp[136]+tmp[14]*tmp[135]+tmp[15]*tmp[134]+tmp[16]*tmp[133]+tmp[17]*tmp[132]+tmp[18]*tmp[131]+tmp[19]*tmp[130]+tmp[20]*tmp[129]+tmp[21]*tmp[128]+tmp[22]*tmp[127]+tmp[23]*tmp[126]+tmp[24]*tmp[125]+tmp[25]*tmp[124]+tmp[26]*tmp[123]+tmp[27]*tmp[122]+tmp[28]*tmp[121]+tmp[29]*tmp[120]+tmp[30]*tmp[119]+tmp[31]*tmp[118]+tmp[32]*tmp[117]+tmp[33]*tmp[116]+tmp[34]*tmp[115]+tmp[35]*tmp[114]+tmp[36]*tmp[113]+tmp[37]*tmp[112]+tmp[38]*tmp[111]+tmp[39]*tmp[110]+tmp[40]*tmp[109]+tmp[41]*tmp[108]+tmp[42]*tmp[107]+tmp[43]*tmp[106]+tmp[44]*tmp[105]+tmp[45]*tmp[104]+tmp[46]*tmp[103]+tmp[47]*tmp[102]+tmp[48]*tmp[101]+tmp[49]*tmp[100];
				ans[50]<=tmp[0]*tmp[150]+tmp[1]*tmp[149]+tmp[2]*tmp[148]+tmp[3]*tmp[147]+tmp[4]*tmp[146]+tmp[5]*tmp[145]+tmp[6]*tmp[144]+tmp[7]*tmp[143]+tmp[8]*tmp[142]+tmp[9]*tmp[141]+tmp[10]*tmp[140]+tmp[11]*tmp[139]+tmp[12]*tmp[138]+tmp[13]*tmp[137]+tmp[14]*tmp[136]+tmp[15]*tmp[135]+tmp[16]*tmp[134]+tmp[17]*tmp[133]+tmp[18]*tmp[132]+tmp[19]*tmp[131]+tmp[20]*tmp[130]+tmp[21]*tmp[129]+tmp[22]*tmp[128]+tmp[23]*tmp[127]+tmp[24]*tmp[126]+tmp[25]*tmp[125]+tmp[26]*tmp[124]+tmp[27]*tmp[123]+tmp[28]*tmp[122]+tmp[29]*tmp[121]+tmp[30]*tmp[120]+tmp[31]*tmp[119]+tmp[32]*tmp[118]+tmp[33]*tmp[117]+tmp[34]*tmp[116]+tmp[35]*tmp[115]+tmp[36]*tmp[114]+tmp[37]*tmp[113]+tmp[38]*tmp[112]+tmp[39]*tmp[111]+tmp[40]*tmp[110]+tmp[41]*tmp[109]+tmp[42]*tmp[108]+tmp[43]*tmp[107]+tmp[44]*tmp[106]+tmp[45]*tmp[105]+tmp[46]*tmp[104]+tmp[47]*tmp[103]+tmp[48]*tmp[102]+tmp[49]*tmp[101]+tmp[50]*tmp[100];
				ans[51]<=tmp[0]*tmp[151]+tmp[1]*tmp[150]+tmp[2]*tmp[149]+tmp[3]*tmp[148]+tmp[4]*tmp[147]+tmp[5]*tmp[146]+tmp[6]*tmp[145]+tmp[7]*tmp[144]+tmp[8]*tmp[143]+tmp[9]*tmp[142]+tmp[10]*tmp[141]+tmp[11]*tmp[140]+tmp[12]*tmp[139]+tmp[13]*tmp[138]+tmp[14]*tmp[137]+tmp[15]*tmp[136]+tmp[16]*tmp[135]+tmp[17]*tmp[134]+tmp[18]*tmp[133]+tmp[19]*tmp[132]+tmp[20]*tmp[131]+tmp[21]*tmp[130]+tmp[22]*tmp[129]+tmp[23]*tmp[128]+tmp[24]*tmp[127]+tmp[25]*tmp[126]+tmp[26]*tmp[125]+tmp[27]*tmp[124]+tmp[28]*tmp[123]+tmp[29]*tmp[122]+tmp[30]*tmp[121]+tmp[31]*tmp[120]+tmp[32]*tmp[119]+tmp[33]*tmp[118]+tmp[34]*tmp[117]+tmp[35]*tmp[116]+tmp[36]*tmp[115]+tmp[37]*tmp[114]+tmp[38]*tmp[113]+tmp[39]*tmp[112]+tmp[40]*tmp[111]+tmp[41]*tmp[110]+tmp[42]*tmp[109]+tmp[43]*tmp[108]+tmp[44]*tmp[107]+tmp[45]*tmp[106]+tmp[46]*tmp[105]+tmp[47]*tmp[104]+tmp[48]*tmp[103]+tmp[49]*tmp[102]+tmp[50]*tmp[101]+tmp[51]*tmp[100];
				ans[52]<=tmp[0]*tmp[152]+tmp[1]*tmp[151]+tmp[2]*tmp[150]+tmp[3]*tmp[149]+tmp[4]*tmp[148]+tmp[5]*tmp[147]+tmp[6]*tmp[146]+tmp[7]*tmp[145]+tmp[8]*tmp[144]+tmp[9]*tmp[143]+tmp[10]*tmp[142]+tmp[11]*tmp[141]+tmp[12]*tmp[140]+tmp[13]*tmp[139]+tmp[14]*tmp[138]+tmp[15]*tmp[137]+tmp[16]*tmp[136]+tmp[17]*tmp[135]+tmp[18]*tmp[134]+tmp[19]*tmp[133]+tmp[20]*tmp[132]+tmp[21]*tmp[131]+tmp[22]*tmp[130]+tmp[23]*tmp[129]+tmp[24]*tmp[128]+tmp[25]*tmp[127]+tmp[26]*tmp[126]+tmp[27]*tmp[125]+tmp[28]*tmp[124]+tmp[29]*tmp[123]+tmp[30]*tmp[122]+tmp[31]*tmp[121]+tmp[32]*tmp[120]+tmp[33]*tmp[119]+tmp[34]*tmp[118]+tmp[35]*tmp[117]+tmp[36]*tmp[116]+tmp[37]*tmp[115]+tmp[38]*tmp[114]+tmp[39]*tmp[113]+tmp[40]*tmp[112]+tmp[41]*tmp[111]+tmp[42]*tmp[110]+tmp[43]*tmp[109]+tmp[44]*tmp[108]+tmp[45]*tmp[107]+tmp[46]*tmp[106]+tmp[47]*tmp[105]+tmp[48]*tmp[104]+tmp[49]*tmp[103]+tmp[50]*tmp[102]+tmp[51]*tmp[101]+tmp[52]*tmp[100];
				ans[53]<=tmp[0]*tmp[153]+tmp[1]*tmp[152]+tmp[2]*tmp[151]+tmp[3]*tmp[150]+tmp[4]*tmp[149]+tmp[5]*tmp[148]+tmp[6]*tmp[147]+tmp[7]*tmp[146]+tmp[8]*tmp[145]+tmp[9]*tmp[144]+tmp[10]*tmp[143]+tmp[11]*tmp[142]+tmp[12]*tmp[141]+tmp[13]*tmp[140]+tmp[14]*tmp[139]+tmp[15]*tmp[138]+tmp[16]*tmp[137]+tmp[17]*tmp[136]+tmp[18]*tmp[135]+tmp[19]*tmp[134]+tmp[20]*tmp[133]+tmp[21]*tmp[132]+tmp[22]*tmp[131]+tmp[23]*tmp[130]+tmp[24]*tmp[129]+tmp[25]*tmp[128]+tmp[26]*tmp[127]+tmp[27]*tmp[126]+tmp[28]*tmp[125]+tmp[29]*tmp[124]+tmp[30]*tmp[123]+tmp[31]*tmp[122]+tmp[32]*tmp[121]+tmp[33]*tmp[120]+tmp[34]*tmp[119]+tmp[35]*tmp[118]+tmp[36]*tmp[117]+tmp[37]*tmp[116]+tmp[38]*tmp[115]+tmp[39]*tmp[114]+tmp[40]*tmp[113]+tmp[41]*tmp[112]+tmp[42]*tmp[111]+tmp[43]*tmp[110]+tmp[44]*tmp[109]+tmp[45]*tmp[108]+tmp[46]*tmp[107]+tmp[47]*tmp[106]+tmp[48]*tmp[105]+tmp[49]*tmp[104]+tmp[50]*tmp[103]+tmp[51]*tmp[102]+tmp[52]*tmp[101]+tmp[53]*tmp[100];
				ans[54]<=tmp[0]*tmp[154]+tmp[1]*tmp[153]+tmp[2]*tmp[152]+tmp[3]*tmp[151]+tmp[4]*tmp[150]+tmp[5]*tmp[149]+tmp[6]*tmp[148]+tmp[7]*tmp[147]+tmp[8]*tmp[146]+tmp[9]*tmp[145]+tmp[10]*tmp[144]+tmp[11]*tmp[143]+tmp[12]*tmp[142]+tmp[13]*tmp[141]+tmp[14]*tmp[140]+tmp[15]*tmp[139]+tmp[16]*tmp[138]+tmp[17]*tmp[137]+tmp[18]*tmp[136]+tmp[19]*tmp[135]+tmp[20]*tmp[134]+tmp[21]*tmp[133]+tmp[22]*tmp[132]+tmp[23]*tmp[131]+tmp[24]*tmp[130]+tmp[25]*tmp[129]+tmp[26]*tmp[128]+tmp[27]*tmp[127]+tmp[28]*tmp[126]+tmp[29]*tmp[125]+tmp[30]*tmp[124]+tmp[31]*tmp[123]+tmp[32]*tmp[122]+tmp[33]*tmp[121]+tmp[34]*tmp[120]+tmp[35]*tmp[119]+tmp[36]*tmp[118]+tmp[37]*tmp[117]+tmp[38]*tmp[116]+tmp[39]*tmp[115]+tmp[40]*tmp[114]+tmp[41]*tmp[113]+tmp[42]*tmp[112]+tmp[43]*tmp[111]+tmp[44]*tmp[110]+tmp[45]*tmp[109]+tmp[46]*tmp[108]+tmp[47]*tmp[107]+tmp[48]*tmp[106]+tmp[49]*tmp[105]+tmp[50]*tmp[104]+tmp[51]*tmp[103]+tmp[52]*tmp[102]+tmp[53]*tmp[101]+tmp[54]*tmp[100];
				ans[55]<=tmp[0]*tmp[155]+tmp[1]*tmp[154]+tmp[2]*tmp[153]+tmp[3]*tmp[152]+tmp[4]*tmp[151]+tmp[5]*tmp[150]+tmp[6]*tmp[149]+tmp[7]*tmp[148]+tmp[8]*tmp[147]+tmp[9]*tmp[146]+tmp[10]*tmp[145]+tmp[11]*tmp[144]+tmp[12]*tmp[143]+tmp[13]*tmp[142]+tmp[14]*tmp[141]+tmp[15]*tmp[140]+tmp[16]*tmp[139]+tmp[17]*tmp[138]+tmp[18]*tmp[137]+tmp[19]*tmp[136]+tmp[20]*tmp[135]+tmp[21]*tmp[134]+tmp[22]*tmp[133]+tmp[23]*tmp[132]+tmp[24]*tmp[131]+tmp[25]*tmp[130]+tmp[26]*tmp[129]+tmp[27]*tmp[128]+tmp[28]*tmp[127]+tmp[29]*tmp[126]+tmp[30]*tmp[125]+tmp[31]*tmp[124]+tmp[32]*tmp[123]+tmp[33]*tmp[122]+tmp[34]*tmp[121]+tmp[35]*tmp[120]+tmp[36]*tmp[119]+tmp[37]*tmp[118]+tmp[38]*tmp[117]+tmp[39]*tmp[116]+tmp[40]*tmp[115]+tmp[41]*tmp[114]+tmp[42]*tmp[113]+tmp[43]*tmp[112]+tmp[44]*tmp[111]+tmp[45]*tmp[110]+tmp[46]*tmp[109]+tmp[47]*tmp[108]+tmp[48]*tmp[107]+tmp[49]*tmp[106]+tmp[50]*tmp[105]+tmp[51]*tmp[104]+tmp[52]*tmp[103]+tmp[53]*tmp[102]+tmp[54]*tmp[101]+tmp[55]*tmp[100];
				ans[56]<=tmp[0]*tmp[156]+tmp[1]*tmp[155]+tmp[2]*tmp[154]+tmp[3]*tmp[153]+tmp[4]*tmp[152]+tmp[5]*tmp[151]+tmp[6]*tmp[150]+tmp[7]*tmp[149]+tmp[8]*tmp[148]+tmp[9]*tmp[147]+tmp[10]*tmp[146]+tmp[11]*tmp[145]+tmp[12]*tmp[144]+tmp[13]*tmp[143]+tmp[14]*tmp[142]+tmp[15]*tmp[141]+tmp[16]*tmp[140]+tmp[17]*tmp[139]+tmp[18]*tmp[138]+tmp[19]*tmp[137]+tmp[20]*tmp[136]+tmp[21]*tmp[135]+tmp[22]*tmp[134]+tmp[23]*tmp[133]+tmp[24]*tmp[132]+tmp[25]*tmp[131]+tmp[26]*tmp[130]+tmp[27]*tmp[129]+tmp[28]*tmp[128]+tmp[29]*tmp[127]+tmp[30]*tmp[126]+tmp[31]*tmp[125]+tmp[32]*tmp[124]+tmp[33]*tmp[123]+tmp[34]*tmp[122]+tmp[35]*tmp[121]+tmp[36]*tmp[120]+tmp[37]*tmp[119]+tmp[38]*tmp[118]+tmp[39]*tmp[117]+tmp[40]*tmp[116]+tmp[41]*tmp[115]+tmp[42]*tmp[114]+tmp[43]*tmp[113]+tmp[44]*tmp[112]+tmp[45]*tmp[111]+tmp[46]*tmp[110]+tmp[47]*tmp[109]+tmp[48]*tmp[108]+tmp[49]*tmp[107]+tmp[50]*tmp[106]+tmp[51]*tmp[105]+tmp[52]*tmp[104]+tmp[53]*tmp[103]+tmp[54]*tmp[102]+tmp[55]*tmp[101]+tmp[56]*tmp[100];
				ans[57]<=tmp[0]*tmp[157]+tmp[1]*tmp[156]+tmp[2]*tmp[155]+tmp[3]*tmp[154]+tmp[4]*tmp[153]+tmp[5]*tmp[152]+tmp[6]*tmp[151]+tmp[7]*tmp[150]+tmp[8]*tmp[149]+tmp[9]*tmp[148]+tmp[10]*tmp[147]+tmp[11]*tmp[146]+tmp[12]*tmp[145]+tmp[13]*tmp[144]+tmp[14]*tmp[143]+tmp[15]*tmp[142]+tmp[16]*tmp[141]+tmp[17]*tmp[140]+tmp[18]*tmp[139]+tmp[19]*tmp[138]+tmp[20]*tmp[137]+tmp[21]*tmp[136]+tmp[22]*tmp[135]+tmp[23]*tmp[134]+tmp[24]*tmp[133]+tmp[25]*tmp[132]+tmp[26]*tmp[131]+tmp[27]*tmp[130]+tmp[28]*tmp[129]+tmp[29]*tmp[128]+tmp[30]*tmp[127]+tmp[31]*tmp[126]+tmp[32]*tmp[125]+tmp[33]*tmp[124]+tmp[34]*tmp[123]+tmp[35]*tmp[122]+tmp[36]*tmp[121]+tmp[37]*tmp[120]+tmp[38]*tmp[119]+tmp[39]*tmp[118]+tmp[40]*tmp[117]+tmp[41]*tmp[116]+tmp[42]*tmp[115]+tmp[43]*tmp[114]+tmp[44]*tmp[113]+tmp[45]*tmp[112]+tmp[46]*tmp[111]+tmp[47]*tmp[110]+tmp[48]*tmp[109]+tmp[49]*tmp[108]+tmp[50]*tmp[107]+tmp[51]*tmp[106]+tmp[52]*tmp[105]+tmp[53]*tmp[104]+tmp[54]*tmp[103]+tmp[55]*tmp[102]+tmp[56]*tmp[101]+tmp[57]*tmp[100];
				ans[58]<=tmp[0]*tmp[158]+tmp[1]*tmp[157]+tmp[2]*tmp[156]+tmp[3]*tmp[155]+tmp[4]*tmp[154]+tmp[5]*tmp[153]+tmp[6]*tmp[152]+tmp[7]*tmp[151]+tmp[8]*tmp[150]+tmp[9]*tmp[149]+tmp[10]*tmp[148]+tmp[11]*tmp[147]+tmp[12]*tmp[146]+tmp[13]*tmp[145]+tmp[14]*tmp[144]+tmp[15]*tmp[143]+tmp[16]*tmp[142]+tmp[17]*tmp[141]+tmp[18]*tmp[140]+tmp[19]*tmp[139]+tmp[20]*tmp[138]+tmp[21]*tmp[137]+tmp[22]*tmp[136]+tmp[23]*tmp[135]+tmp[24]*tmp[134]+tmp[25]*tmp[133]+tmp[26]*tmp[132]+tmp[27]*tmp[131]+tmp[28]*tmp[130]+tmp[29]*tmp[129]+tmp[30]*tmp[128]+tmp[31]*tmp[127]+tmp[32]*tmp[126]+tmp[33]*tmp[125]+tmp[34]*tmp[124]+tmp[35]*tmp[123]+tmp[36]*tmp[122]+tmp[37]*tmp[121]+tmp[38]*tmp[120]+tmp[39]*tmp[119]+tmp[40]*tmp[118]+tmp[41]*tmp[117]+tmp[42]*tmp[116]+tmp[43]*tmp[115]+tmp[44]*tmp[114]+tmp[45]*tmp[113]+tmp[46]*tmp[112]+tmp[47]*tmp[111]+tmp[48]*tmp[110]+tmp[49]*tmp[109]+tmp[50]*tmp[108]+tmp[51]*tmp[107]+tmp[52]*tmp[106]+tmp[53]*tmp[105]+tmp[54]*tmp[104]+tmp[55]*tmp[103]+tmp[56]*tmp[102]+tmp[57]*tmp[101]+tmp[58]*tmp[100];
				ans[59]<=tmp[0]*tmp[159]+tmp[1]*tmp[158]+tmp[2]*tmp[157]+tmp[3]*tmp[156]+tmp[4]*tmp[155]+tmp[5]*tmp[154]+tmp[6]*tmp[153]+tmp[7]*tmp[152]+tmp[8]*tmp[151]+tmp[9]*tmp[150]+tmp[10]*tmp[149]+tmp[11]*tmp[148]+tmp[12]*tmp[147]+tmp[13]*tmp[146]+tmp[14]*tmp[145]+tmp[15]*tmp[144]+tmp[16]*tmp[143]+tmp[17]*tmp[142]+tmp[18]*tmp[141]+tmp[19]*tmp[140]+tmp[20]*tmp[139]+tmp[21]*tmp[138]+tmp[22]*tmp[137]+tmp[23]*tmp[136]+tmp[24]*tmp[135]+tmp[25]*tmp[134]+tmp[26]*tmp[133]+tmp[27]*tmp[132]+tmp[28]*tmp[131]+tmp[29]*tmp[130]+tmp[30]*tmp[129]+tmp[31]*tmp[128]+tmp[32]*tmp[127]+tmp[33]*tmp[126]+tmp[34]*tmp[125]+tmp[35]*tmp[124]+tmp[36]*tmp[123]+tmp[37]*tmp[122]+tmp[38]*tmp[121]+tmp[39]*tmp[120]+tmp[40]*tmp[119]+tmp[41]*tmp[118]+tmp[42]*tmp[117]+tmp[43]*tmp[116]+tmp[44]*tmp[115]+tmp[45]*tmp[114]+tmp[46]*tmp[113]+tmp[47]*tmp[112]+tmp[48]*tmp[111]+tmp[49]*tmp[110]+tmp[50]*tmp[109]+tmp[51]*tmp[108]+tmp[52]*tmp[107]+tmp[53]*tmp[106]+tmp[54]*tmp[105]+tmp[55]*tmp[104]+tmp[56]*tmp[103]+tmp[57]*tmp[102]+tmp[58]*tmp[101]+tmp[59]*tmp[100];
				ans[60]<=tmp[0]*tmp[160]+tmp[1]*tmp[159]+tmp[2]*tmp[158]+tmp[3]*tmp[157]+tmp[4]*tmp[156]+tmp[5]*tmp[155]+tmp[6]*tmp[154]+tmp[7]*tmp[153]+tmp[8]*tmp[152]+tmp[9]*tmp[151]+tmp[10]*tmp[150]+tmp[11]*tmp[149]+tmp[12]*tmp[148]+tmp[13]*tmp[147]+tmp[14]*tmp[146]+tmp[15]*tmp[145]+tmp[16]*tmp[144]+tmp[17]*tmp[143]+tmp[18]*tmp[142]+tmp[19]*tmp[141]+tmp[20]*tmp[140]+tmp[21]*tmp[139]+tmp[22]*tmp[138]+tmp[23]*tmp[137]+tmp[24]*tmp[136]+tmp[25]*tmp[135]+tmp[26]*tmp[134]+tmp[27]*tmp[133]+tmp[28]*tmp[132]+tmp[29]*tmp[131]+tmp[30]*tmp[130]+tmp[31]*tmp[129]+tmp[32]*tmp[128]+tmp[33]*tmp[127]+tmp[34]*tmp[126]+tmp[35]*tmp[125]+tmp[36]*tmp[124]+tmp[37]*tmp[123]+tmp[38]*tmp[122]+tmp[39]*tmp[121]+tmp[40]*tmp[120]+tmp[41]*tmp[119]+tmp[42]*tmp[118]+tmp[43]*tmp[117]+tmp[44]*tmp[116]+tmp[45]*tmp[115]+tmp[46]*tmp[114]+tmp[47]*tmp[113]+tmp[48]*tmp[112]+tmp[49]*tmp[111]+tmp[50]*tmp[110]+tmp[51]*tmp[109]+tmp[52]*tmp[108]+tmp[53]*tmp[107]+tmp[54]*tmp[106]+tmp[55]*tmp[105]+tmp[56]*tmp[104]+tmp[57]*tmp[103]+tmp[58]*tmp[102]+tmp[59]*tmp[101]+tmp[60]*tmp[100];
				ans[61]<=tmp[0]*tmp[161]+tmp[1]*tmp[160]+tmp[2]*tmp[159]+tmp[3]*tmp[158]+tmp[4]*tmp[157]+tmp[5]*tmp[156]+tmp[6]*tmp[155]+tmp[7]*tmp[154]+tmp[8]*tmp[153]+tmp[9]*tmp[152]+tmp[10]*tmp[151]+tmp[11]*tmp[150]+tmp[12]*tmp[149]+tmp[13]*tmp[148]+tmp[14]*tmp[147]+tmp[15]*tmp[146]+tmp[16]*tmp[145]+tmp[17]*tmp[144]+tmp[18]*tmp[143]+tmp[19]*tmp[142]+tmp[20]*tmp[141]+tmp[21]*tmp[140]+tmp[22]*tmp[139]+tmp[23]*tmp[138]+tmp[24]*tmp[137]+tmp[25]*tmp[136]+tmp[26]*tmp[135]+tmp[27]*tmp[134]+tmp[28]*tmp[133]+tmp[29]*tmp[132]+tmp[30]*tmp[131]+tmp[31]*tmp[130]+tmp[32]*tmp[129]+tmp[33]*tmp[128]+tmp[34]*tmp[127]+tmp[35]*tmp[126]+tmp[36]*tmp[125]+tmp[37]*tmp[124]+tmp[38]*tmp[123]+tmp[39]*tmp[122]+tmp[40]*tmp[121]+tmp[41]*tmp[120]+tmp[42]*tmp[119]+tmp[43]*tmp[118]+tmp[44]*tmp[117]+tmp[45]*tmp[116]+tmp[46]*tmp[115]+tmp[47]*tmp[114]+tmp[48]*tmp[113]+tmp[49]*tmp[112]+tmp[50]*tmp[111]+tmp[51]*tmp[110]+tmp[52]*tmp[109]+tmp[53]*tmp[108]+tmp[54]*tmp[107]+tmp[55]*tmp[106]+tmp[56]*tmp[105]+tmp[57]*tmp[104]+tmp[58]*tmp[103]+tmp[59]*tmp[102]+tmp[60]*tmp[101]+tmp[61]*tmp[100];
				ans[62]<=tmp[0]*tmp[162]+tmp[1]*tmp[161]+tmp[2]*tmp[160]+tmp[3]*tmp[159]+tmp[4]*tmp[158]+tmp[5]*tmp[157]+tmp[6]*tmp[156]+tmp[7]*tmp[155]+tmp[8]*tmp[154]+tmp[9]*tmp[153]+tmp[10]*tmp[152]+tmp[11]*tmp[151]+tmp[12]*tmp[150]+tmp[13]*tmp[149]+tmp[14]*tmp[148]+tmp[15]*tmp[147]+tmp[16]*tmp[146]+tmp[17]*tmp[145]+tmp[18]*tmp[144]+tmp[19]*tmp[143]+tmp[20]*tmp[142]+tmp[21]*tmp[141]+tmp[22]*tmp[140]+tmp[23]*tmp[139]+tmp[24]*tmp[138]+tmp[25]*tmp[137]+tmp[26]*tmp[136]+tmp[27]*tmp[135]+tmp[28]*tmp[134]+tmp[29]*tmp[133]+tmp[30]*tmp[132]+tmp[31]*tmp[131]+tmp[32]*tmp[130]+tmp[33]*tmp[129]+tmp[34]*tmp[128]+tmp[35]*tmp[127]+tmp[36]*tmp[126]+tmp[37]*tmp[125]+tmp[38]*tmp[124]+tmp[39]*tmp[123]+tmp[40]*tmp[122]+tmp[41]*tmp[121]+tmp[42]*tmp[120]+tmp[43]*tmp[119]+tmp[44]*tmp[118]+tmp[45]*tmp[117]+tmp[46]*tmp[116]+tmp[47]*tmp[115]+tmp[48]*tmp[114]+tmp[49]*tmp[113]+tmp[50]*tmp[112]+tmp[51]*tmp[111]+tmp[52]*tmp[110]+tmp[53]*tmp[109]+tmp[54]*tmp[108]+tmp[55]*tmp[107]+tmp[56]*tmp[106]+tmp[57]*tmp[105]+tmp[58]*tmp[104]+tmp[59]*tmp[103]+tmp[60]*tmp[102]+tmp[61]*tmp[101]+tmp[62]*tmp[100];
				ans[63]<=tmp[0]*tmp[163]+tmp[1]*tmp[162]+tmp[2]*tmp[161]+tmp[3]*tmp[160]+tmp[4]*tmp[159]+tmp[5]*tmp[158]+tmp[6]*tmp[157]+tmp[7]*tmp[156]+tmp[8]*tmp[155]+tmp[9]*tmp[154]+tmp[10]*tmp[153]+tmp[11]*tmp[152]+tmp[12]*tmp[151]+tmp[13]*tmp[150]+tmp[14]*tmp[149]+tmp[15]*tmp[148]+tmp[16]*tmp[147]+tmp[17]*tmp[146]+tmp[18]*tmp[145]+tmp[19]*tmp[144]+tmp[20]*tmp[143]+tmp[21]*tmp[142]+tmp[22]*tmp[141]+tmp[23]*tmp[140]+tmp[24]*tmp[139]+tmp[25]*tmp[138]+tmp[26]*tmp[137]+tmp[27]*tmp[136]+tmp[28]*tmp[135]+tmp[29]*tmp[134]+tmp[30]*tmp[133]+tmp[31]*tmp[132]+tmp[32]*tmp[131]+tmp[33]*tmp[130]+tmp[34]*tmp[129]+tmp[35]*tmp[128]+tmp[36]*tmp[127]+tmp[37]*tmp[126]+tmp[38]*tmp[125]+tmp[39]*tmp[124]+tmp[40]*tmp[123]+tmp[41]*tmp[122]+tmp[42]*tmp[121]+tmp[43]*tmp[120]+tmp[44]*tmp[119]+tmp[45]*tmp[118]+tmp[46]*tmp[117]+tmp[47]*tmp[116]+tmp[48]*tmp[115]+tmp[49]*tmp[114]+tmp[50]*tmp[113]+tmp[51]*tmp[112]+tmp[52]*tmp[111]+tmp[53]*tmp[110]+tmp[54]*tmp[109]+tmp[55]*tmp[108]+tmp[56]*tmp[107]+tmp[57]*tmp[106]+tmp[58]*tmp[105]+tmp[59]*tmp[104]+tmp[60]*tmp[103]+tmp[61]*tmp[102]+tmp[62]*tmp[101]+tmp[63]*tmp[100];
				ans[64]<=tmp[0]*tmp[164]+tmp[1]*tmp[163]+tmp[2]*tmp[162]+tmp[3]*tmp[161]+tmp[4]*tmp[160]+tmp[5]*tmp[159]+tmp[6]*tmp[158]+tmp[7]*tmp[157]+tmp[8]*tmp[156]+tmp[9]*tmp[155]+tmp[10]*tmp[154]+tmp[11]*tmp[153]+tmp[12]*tmp[152]+tmp[13]*tmp[151]+tmp[14]*tmp[150]+tmp[15]*tmp[149]+tmp[16]*tmp[148]+tmp[17]*tmp[147]+tmp[18]*tmp[146]+tmp[19]*tmp[145]+tmp[20]*tmp[144]+tmp[21]*tmp[143]+tmp[22]*tmp[142]+tmp[23]*tmp[141]+tmp[24]*tmp[140]+tmp[25]*tmp[139]+tmp[26]*tmp[138]+tmp[27]*tmp[137]+tmp[28]*tmp[136]+tmp[29]*tmp[135]+tmp[30]*tmp[134]+tmp[31]*tmp[133]+tmp[32]*tmp[132]+tmp[33]*tmp[131]+tmp[34]*tmp[130]+tmp[35]*tmp[129]+tmp[36]*tmp[128]+tmp[37]*tmp[127]+tmp[38]*tmp[126]+tmp[39]*tmp[125]+tmp[40]*tmp[124]+tmp[41]*tmp[123]+tmp[42]*tmp[122]+tmp[43]*tmp[121]+tmp[44]*tmp[120]+tmp[45]*tmp[119]+tmp[46]*tmp[118]+tmp[47]*tmp[117]+tmp[48]*tmp[116]+tmp[49]*tmp[115]+tmp[50]*tmp[114]+tmp[51]*tmp[113]+tmp[52]*tmp[112]+tmp[53]*tmp[111]+tmp[54]*tmp[110]+tmp[55]*tmp[109]+tmp[56]*tmp[108]+tmp[57]*tmp[107]+tmp[58]*tmp[106]+tmp[59]*tmp[105]+tmp[60]*tmp[104]+tmp[61]*tmp[103]+tmp[62]*tmp[102]+tmp[63]*tmp[101]+tmp[64]*tmp[100];
				ans[65]<=tmp[0]*tmp[165]+tmp[1]*tmp[164]+tmp[2]*tmp[163]+tmp[3]*tmp[162]+tmp[4]*tmp[161]+tmp[5]*tmp[160]+tmp[6]*tmp[159]+tmp[7]*tmp[158]+tmp[8]*tmp[157]+tmp[9]*tmp[156]+tmp[10]*tmp[155]+tmp[11]*tmp[154]+tmp[12]*tmp[153]+tmp[13]*tmp[152]+tmp[14]*tmp[151]+tmp[15]*tmp[150]+tmp[16]*tmp[149]+tmp[17]*tmp[148]+tmp[18]*tmp[147]+tmp[19]*tmp[146]+tmp[20]*tmp[145]+tmp[21]*tmp[144]+tmp[22]*tmp[143]+tmp[23]*tmp[142]+tmp[24]*tmp[141]+tmp[25]*tmp[140]+tmp[26]*tmp[139]+tmp[27]*tmp[138]+tmp[28]*tmp[137]+tmp[29]*tmp[136]+tmp[30]*tmp[135]+tmp[31]*tmp[134]+tmp[32]*tmp[133]+tmp[33]*tmp[132]+tmp[34]*tmp[131]+tmp[35]*tmp[130]+tmp[36]*tmp[129]+tmp[37]*tmp[128]+tmp[38]*tmp[127]+tmp[39]*tmp[126]+tmp[40]*tmp[125]+tmp[41]*tmp[124]+tmp[42]*tmp[123]+tmp[43]*tmp[122]+tmp[44]*tmp[121]+tmp[45]*tmp[120]+tmp[46]*tmp[119]+tmp[47]*tmp[118]+tmp[48]*tmp[117]+tmp[49]*tmp[116]+tmp[50]*tmp[115]+tmp[51]*tmp[114]+tmp[52]*tmp[113]+tmp[53]*tmp[112]+tmp[54]*tmp[111]+tmp[55]*tmp[110]+tmp[56]*tmp[109]+tmp[57]*tmp[108]+tmp[58]*tmp[107]+tmp[59]*tmp[106]+tmp[60]*tmp[105]+tmp[61]*tmp[104]+tmp[62]*tmp[103]+tmp[63]*tmp[102]+tmp[64]*tmp[101]+tmp[65]*tmp[100];
				ans[66]<=tmp[0]*tmp[166]+tmp[1]*tmp[165]+tmp[2]*tmp[164]+tmp[3]*tmp[163]+tmp[4]*tmp[162]+tmp[5]*tmp[161]+tmp[6]*tmp[160]+tmp[7]*tmp[159]+tmp[8]*tmp[158]+tmp[9]*tmp[157]+tmp[10]*tmp[156]+tmp[11]*tmp[155]+tmp[12]*tmp[154]+tmp[13]*tmp[153]+tmp[14]*tmp[152]+tmp[15]*tmp[151]+tmp[16]*tmp[150]+tmp[17]*tmp[149]+tmp[18]*tmp[148]+tmp[19]*tmp[147]+tmp[20]*tmp[146]+tmp[21]*tmp[145]+tmp[22]*tmp[144]+tmp[23]*tmp[143]+tmp[24]*tmp[142]+tmp[25]*tmp[141]+tmp[26]*tmp[140]+tmp[27]*tmp[139]+tmp[28]*tmp[138]+tmp[29]*tmp[137]+tmp[30]*tmp[136]+tmp[31]*tmp[135]+tmp[32]*tmp[134]+tmp[33]*tmp[133]+tmp[34]*tmp[132]+tmp[35]*tmp[131]+tmp[36]*tmp[130]+tmp[37]*tmp[129]+tmp[38]*tmp[128]+tmp[39]*tmp[127]+tmp[40]*tmp[126]+tmp[41]*tmp[125]+tmp[42]*tmp[124]+tmp[43]*tmp[123]+tmp[44]*tmp[122]+tmp[45]*tmp[121]+tmp[46]*tmp[120]+tmp[47]*tmp[119]+tmp[48]*tmp[118]+tmp[49]*tmp[117]+tmp[50]*tmp[116]+tmp[51]*tmp[115]+tmp[52]*tmp[114]+tmp[53]*tmp[113]+tmp[54]*tmp[112]+tmp[55]*tmp[111]+tmp[56]*tmp[110]+tmp[57]*tmp[109]+tmp[58]*tmp[108]+tmp[59]*tmp[107]+tmp[60]*tmp[106]+tmp[61]*tmp[105]+tmp[62]*tmp[104]+tmp[63]*tmp[103]+tmp[64]*tmp[102]+tmp[65]*tmp[101]+tmp[66]*tmp[100];
				ans[67]<=tmp[0]*tmp[167]+tmp[1]*tmp[166]+tmp[2]*tmp[165]+tmp[3]*tmp[164]+tmp[4]*tmp[163]+tmp[5]*tmp[162]+tmp[6]*tmp[161]+tmp[7]*tmp[160]+tmp[8]*tmp[159]+tmp[9]*tmp[158]+tmp[10]*tmp[157]+tmp[11]*tmp[156]+tmp[12]*tmp[155]+tmp[13]*tmp[154]+tmp[14]*tmp[153]+tmp[15]*tmp[152]+tmp[16]*tmp[151]+tmp[17]*tmp[150]+tmp[18]*tmp[149]+tmp[19]*tmp[148]+tmp[20]*tmp[147]+tmp[21]*tmp[146]+tmp[22]*tmp[145]+tmp[23]*tmp[144]+tmp[24]*tmp[143]+tmp[25]*tmp[142]+tmp[26]*tmp[141]+tmp[27]*tmp[140]+tmp[28]*tmp[139]+tmp[29]*tmp[138]+tmp[30]*tmp[137]+tmp[31]*tmp[136]+tmp[32]*tmp[135]+tmp[33]*tmp[134]+tmp[34]*tmp[133]+tmp[35]*tmp[132]+tmp[36]*tmp[131]+tmp[37]*tmp[130]+tmp[38]*tmp[129]+tmp[39]*tmp[128]+tmp[40]*tmp[127]+tmp[41]*tmp[126]+tmp[42]*tmp[125]+tmp[43]*tmp[124]+tmp[44]*tmp[123]+tmp[45]*tmp[122]+tmp[46]*tmp[121]+tmp[47]*tmp[120]+tmp[48]*tmp[119]+tmp[49]*tmp[118]+tmp[50]*tmp[117]+tmp[51]*tmp[116]+tmp[52]*tmp[115]+tmp[53]*tmp[114]+tmp[54]*tmp[113]+tmp[55]*tmp[112]+tmp[56]*tmp[111]+tmp[57]*tmp[110]+tmp[58]*tmp[109]+tmp[59]*tmp[108]+tmp[60]*tmp[107]+tmp[61]*tmp[106]+tmp[62]*tmp[105]+tmp[63]*tmp[104]+tmp[64]*tmp[103]+tmp[65]*tmp[102]+tmp[66]*tmp[101]+tmp[67]*tmp[100];
				ans[68]<=tmp[0]*tmp[168]+tmp[1]*tmp[167]+tmp[2]*tmp[166]+tmp[3]*tmp[165]+tmp[4]*tmp[164]+tmp[5]*tmp[163]+tmp[6]*tmp[162]+tmp[7]*tmp[161]+tmp[8]*tmp[160]+tmp[9]*tmp[159]+tmp[10]*tmp[158]+tmp[11]*tmp[157]+tmp[12]*tmp[156]+tmp[13]*tmp[155]+tmp[14]*tmp[154]+tmp[15]*tmp[153]+tmp[16]*tmp[152]+tmp[17]*tmp[151]+tmp[18]*tmp[150]+tmp[19]*tmp[149]+tmp[20]*tmp[148]+tmp[21]*tmp[147]+tmp[22]*tmp[146]+tmp[23]*tmp[145]+tmp[24]*tmp[144]+tmp[25]*tmp[143]+tmp[26]*tmp[142]+tmp[27]*tmp[141]+tmp[28]*tmp[140]+tmp[29]*tmp[139]+tmp[30]*tmp[138]+tmp[31]*tmp[137]+tmp[32]*tmp[136]+tmp[33]*tmp[135]+tmp[34]*tmp[134]+tmp[35]*tmp[133]+tmp[36]*tmp[132]+tmp[37]*tmp[131]+tmp[38]*tmp[130]+tmp[39]*tmp[129]+tmp[40]*tmp[128]+tmp[41]*tmp[127]+tmp[42]*tmp[126]+tmp[43]*tmp[125]+tmp[44]*tmp[124]+tmp[45]*tmp[123]+tmp[46]*tmp[122]+tmp[47]*tmp[121]+tmp[48]*tmp[120]+tmp[49]*tmp[119]+tmp[50]*tmp[118]+tmp[51]*tmp[117]+tmp[52]*tmp[116]+tmp[53]*tmp[115]+tmp[54]*tmp[114]+tmp[55]*tmp[113]+tmp[56]*tmp[112]+tmp[57]*tmp[111]+tmp[58]*tmp[110]+tmp[59]*tmp[109]+tmp[60]*tmp[108]+tmp[61]*tmp[107]+tmp[62]*tmp[106]+tmp[63]*tmp[105]+tmp[64]*tmp[104]+tmp[65]*tmp[103]+tmp[66]*tmp[102]+tmp[67]*tmp[101]+tmp[68]*tmp[100];
				ans[69]<=tmp[0]*tmp[169]+tmp[1]*tmp[168]+tmp[2]*tmp[167]+tmp[3]*tmp[166]+tmp[4]*tmp[165]+tmp[5]*tmp[164]+tmp[6]*tmp[163]+tmp[7]*tmp[162]+tmp[8]*tmp[161]+tmp[9]*tmp[160]+tmp[10]*tmp[159]+tmp[11]*tmp[158]+tmp[12]*tmp[157]+tmp[13]*tmp[156]+tmp[14]*tmp[155]+tmp[15]*tmp[154]+tmp[16]*tmp[153]+tmp[17]*tmp[152]+tmp[18]*tmp[151]+tmp[19]*tmp[150]+tmp[20]*tmp[149]+tmp[21]*tmp[148]+tmp[22]*tmp[147]+tmp[23]*tmp[146]+tmp[24]*tmp[145]+tmp[25]*tmp[144]+tmp[26]*tmp[143]+tmp[27]*tmp[142]+tmp[28]*tmp[141]+tmp[29]*tmp[140]+tmp[30]*tmp[139]+tmp[31]*tmp[138]+tmp[32]*tmp[137]+tmp[33]*tmp[136]+tmp[34]*tmp[135]+tmp[35]*tmp[134]+tmp[36]*tmp[133]+tmp[37]*tmp[132]+tmp[38]*tmp[131]+tmp[39]*tmp[130]+tmp[40]*tmp[129]+tmp[41]*tmp[128]+tmp[42]*tmp[127]+tmp[43]*tmp[126]+tmp[44]*tmp[125]+tmp[45]*tmp[124]+tmp[46]*tmp[123]+tmp[47]*tmp[122]+tmp[48]*tmp[121]+tmp[49]*tmp[120]+tmp[50]*tmp[119]+tmp[51]*tmp[118]+tmp[52]*tmp[117]+tmp[53]*tmp[116]+tmp[54]*tmp[115]+tmp[55]*tmp[114]+tmp[56]*tmp[113]+tmp[57]*tmp[112]+tmp[58]*tmp[111]+tmp[59]*tmp[110]+tmp[60]*tmp[109]+tmp[61]*tmp[108]+tmp[62]*tmp[107]+tmp[63]*tmp[106]+tmp[64]*tmp[105]+tmp[65]*tmp[104]+tmp[66]*tmp[103]+tmp[67]*tmp[102]+tmp[68]*tmp[101]+tmp[69]*tmp[100];
				ans[70]<=tmp[0]*tmp[170]+tmp[1]*tmp[169]+tmp[2]*tmp[168]+tmp[3]*tmp[167]+tmp[4]*tmp[166]+tmp[5]*tmp[165]+tmp[6]*tmp[164]+tmp[7]*tmp[163]+tmp[8]*tmp[162]+tmp[9]*tmp[161]+tmp[10]*tmp[160]+tmp[11]*tmp[159]+tmp[12]*tmp[158]+tmp[13]*tmp[157]+tmp[14]*tmp[156]+tmp[15]*tmp[155]+tmp[16]*tmp[154]+tmp[17]*tmp[153]+tmp[18]*tmp[152]+tmp[19]*tmp[151]+tmp[20]*tmp[150]+tmp[21]*tmp[149]+tmp[22]*tmp[148]+tmp[23]*tmp[147]+tmp[24]*tmp[146]+tmp[25]*tmp[145]+tmp[26]*tmp[144]+tmp[27]*tmp[143]+tmp[28]*tmp[142]+tmp[29]*tmp[141]+tmp[30]*tmp[140]+tmp[31]*tmp[139]+tmp[32]*tmp[138]+tmp[33]*tmp[137]+tmp[34]*tmp[136]+tmp[35]*tmp[135]+tmp[36]*tmp[134]+tmp[37]*tmp[133]+tmp[38]*tmp[132]+tmp[39]*tmp[131]+tmp[40]*tmp[130]+tmp[41]*tmp[129]+tmp[42]*tmp[128]+tmp[43]*tmp[127]+tmp[44]*tmp[126]+tmp[45]*tmp[125]+tmp[46]*tmp[124]+tmp[47]*tmp[123]+tmp[48]*tmp[122]+tmp[49]*tmp[121]+tmp[50]*tmp[120]+tmp[51]*tmp[119]+tmp[52]*tmp[118]+tmp[53]*tmp[117]+tmp[54]*tmp[116]+tmp[55]*tmp[115]+tmp[56]*tmp[114]+tmp[57]*tmp[113]+tmp[58]*tmp[112]+tmp[59]*tmp[111]+tmp[60]*tmp[110]+tmp[61]*tmp[109]+tmp[62]*tmp[108]+tmp[63]*tmp[107]+tmp[64]*tmp[106]+tmp[65]*tmp[105]+tmp[66]*tmp[104]+tmp[67]*tmp[103]+tmp[68]*tmp[102]+tmp[69]*tmp[101]+tmp[70]*tmp[100];
				ans[71]<=tmp[0]*tmp[171]+tmp[1]*tmp[170]+tmp[2]*tmp[169]+tmp[3]*tmp[168]+tmp[4]*tmp[167]+tmp[5]*tmp[166]+tmp[6]*tmp[165]+tmp[7]*tmp[164]+tmp[8]*tmp[163]+tmp[9]*tmp[162]+tmp[10]*tmp[161]+tmp[11]*tmp[160]+tmp[12]*tmp[159]+tmp[13]*tmp[158]+tmp[14]*tmp[157]+tmp[15]*tmp[156]+tmp[16]*tmp[155]+tmp[17]*tmp[154]+tmp[18]*tmp[153]+tmp[19]*tmp[152]+tmp[20]*tmp[151]+tmp[21]*tmp[150]+tmp[22]*tmp[149]+tmp[23]*tmp[148]+tmp[24]*tmp[147]+tmp[25]*tmp[146]+tmp[26]*tmp[145]+tmp[27]*tmp[144]+tmp[28]*tmp[143]+tmp[29]*tmp[142]+tmp[30]*tmp[141]+tmp[31]*tmp[140]+tmp[32]*tmp[139]+tmp[33]*tmp[138]+tmp[34]*tmp[137]+tmp[35]*tmp[136]+tmp[36]*tmp[135]+tmp[37]*tmp[134]+tmp[38]*tmp[133]+tmp[39]*tmp[132]+tmp[40]*tmp[131]+tmp[41]*tmp[130]+tmp[42]*tmp[129]+tmp[43]*tmp[128]+tmp[44]*tmp[127]+tmp[45]*tmp[126]+tmp[46]*tmp[125]+tmp[47]*tmp[124]+tmp[48]*tmp[123]+tmp[49]*tmp[122]+tmp[50]*tmp[121]+tmp[51]*tmp[120]+tmp[52]*tmp[119]+tmp[53]*tmp[118]+tmp[54]*tmp[117]+tmp[55]*tmp[116]+tmp[56]*tmp[115]+tmp[57]*tmp[114]+tmp[58]*tmp[113]+tmp[59]*tmp[112]+tmp[60]*tmp[111]+tmp[61]*tmp[110]+tmp[62]*tmp[109]+tmp[63]*tmp[108]+tmp[64]*tmp[107]+tmp[65]*tmp[106]+tmp[66]*tmp[105]+tmp[67]*tmp[104]+tmp[68]*tmp[103]+tmp[69]*tmp[102]+tmp[70]*tmp[101]+tmp[71]*tmp[100];
				ans[72]<=tmp[0]*tmp[172]+tmp[1]*tmp[171]+tmp[2]*tmp[170]+tmp[3]*tmp[169]+tmp[4]*tmp[168]+tmp[5]*tmp[167]+tmp[6]*tmp[166]+tmp[7]*tmp[165]+tmp[8]*tmp[164]+tmp[9]*tmp[163]+tmp[10]*tmp[162]+tmp[11]*tmp[161]+tmp[12]*tmp[160]+tmp[13]*tmp[159]+tmp[14]*tmp[158]+tmp[15]*tmp[157]+tmp[16]*tmp[156]+tmp[17]*tmp[155]+tmp[18]*tmp[154]+tmp[19]*tmp[153]+tmp[20]*tmp[152]+tmp[21]*tmp[151]+tmp[22]*tmp[150]+tmp[23]*tmp[149]+tmp[24]*tmp[148]+tmp[25]*tmp[147]+tmp[26]*tmp[146]+tmp[27]*tmp[145]+tmp[28]*tmp[144]+tmp[29]*tmp[143]+tmp[30]*tmp[142]+tmp[31]*tmp[141]+tmp[32]*tmp[140]+tmp[33]*tmp[139]+tmp[34]*tmp[138]+tmp[35]*tmp[137]+tmp[36]*tmp[136]+tmp[37]*tmp[135]+tmp[38]*tmp[134]+tmp[39]*tmp[133]+tmp[40]*tmp[132]+tmp[41]*tmp[131]+tmp[42]*tmp[130]+tmp[43]*tmp[129]+tmp[44]*tmp[128]+tmp[45]*tmp[127]+tmp[46]*tmp[126]+tmp[47]*tmp[125]+tmp[48]*tmp[124]+tmp[49]*tmp[123]+tmp[50]*tmp[122]+tmp[51]*tmp[121]+tmp[52]*tmp[120]+tmp[53]*tmp[119]+tmp[54]*tmp[118]+tmp[55]*tmp[117]+tmp[56]*tmp[116]+tmp[57]*tmp[115]+tmp[58]*tmp[114]+tmp[59]*tmp[113]+tmp[60]*tmp[112]+tmp[61]*tmp[111]+tmp[62]*tmp[110]+tmp[63]*tmp[109]+tmp[64]*tmp[108]+tmp[65]*tmp[107]+tmp[66]*tmp[106]+tmp[67]*tmp[105]+tmp[68]*tmp[104]+tmp[69]*tmp[103]+tmp[70]*tmp[102]+tmp[71]*tmp[101]+tmp[72]*tmp[100];
				ans[73]<=tmp[0]*tmp[173]+tmp[1]*tmp[172]+tmp[2]*tmp[171]+tmp[3]*tmp[170]+tmp[4]*tmp[169]+tmp[5]*tmp[168]+tmp[6]*tmp[167]+tmp[7]*tmp[166]+tmp[8]*tmp[165]+tmp[9]*tmp[164]+tmp[10]*tmp[163]+tmp[11]*tmp[162]+tmp[12]*tmp[161]+tmp[13]*tmp[160]+tmp[14]*tmp[159]+tmp[15]*tmp[158]+tmp[16]*tmp[157]+tmp[17]*tmp[156]+tmp[18]*tmp[155]+tmp[19]*tmp[154]+tmp[20]*tmp[153]+tmp[21]*tmp[152]+tmp[22]*tmp[151]+tmp[23]*tmp[150]+tmp[24]*tmp[149]+tmp[25]*tmp[148]+tmp[26]*tmp[147]+tmp[27]*tmp[146]+tmp[28]*tmp[145]+tmp[29]*tmp[144]+tmp[30]*tmp[143]+tmp[31]*tmp[142]+tmp[32]*tmp[141]+tmp[33]*tmp[140]+tmp[34]*tmp[139]+tmp[35]*tmp[138]+tmp[36]*tmp[137]+tmp[37]*tmp[136]+tmp[38]*tmp[135]+tmp[39]*tmp[134]+tmp[40]*tmp[133]+tmp[41]*tmp[132]+tmp[42]*tmp[131]+tmp[43]*tmp[130]+tmp[44]*tmp[129]+tmp[45]*tmp[128]+tmp[46]*tmp[127]+tmp[47]*tmp[126]+tmp[48]*tmp[125]+tmp[49]*tmp[124]+tmp[50]*tmp[123]+tmp[51]*tmp[122]+tmp[52]*tmp[121]+tmp[53]*tmp[120]+tmp[54]*tmp[119]+tmp[55]*tmp[118]+tmp[56]*tmp[117]+tmp[57]*tmp[116]+tmp[58]*tmp[115]+tmp[59]*tmp[114]+tmp[60]*tmp[113]+tmp[61]*tmp[112]+tmp[62]*tmp[111]+tmp[63]*tmp[110]+tmp[64]*tmp[109]+tmp[65]*tmp[108]+tmp[66]*tmp[107]+tmp[67]*tmp[106]+tmp[68]*tmp[105]+tmp[69]*tmp[104]+tmp[70]*tmp[103]+tmp[71]*tmp[102]+tmp[72]*tmp[101]+tmp[73]*tmp[100];
				ans[74]<=tmp[0]*tmp[174]+tmp[1]*tmp[173]+tmp[2]*tmp[172]+tmp[3]*tmp[171]+tmp[4]*tmp[170]+tmp[5]*tmp[169]+tmp[6]*tmp[168]+tmp[7]*tmp[167]+tmp[8]*tmp[166]+tmp[9]*tmp[165]+tmp[10]*tmp[164]+tmp[11]*tmp[163]+tmp[12]*tmp[162]+tmp[13]*tmp[161]+tmp[14]*tmp[160]+tmp[15]*tmp[159]+tmp[16]*tmp[158]+tmp[17]*tmp[157]+tmp[18]*tmp[156]+tmp[19]*tmp[155]+tmp[20]*tmp[154]+tmp[21]*tmp[153]+tmp[22]*tmp[152]+tmp[23]*tmp[151]+tmp[24]*tmp[150]+tmp[25]*tmp[149]+tmp[26]*tmp[148]+tmp[27]*tmp[147]+tmp[28]*tmp[146]+tmp[29]*tmp[145]+tmp[30]*tmp[144]+tmp[31]*tmp[143]+tmp[32]*tmp[142]+tmp[33]*tmp[141]+tmp[34]*tmp[140]+tmp[35]*tmp[139]+tmp[36]*tmp[138]+tmp[37]*tmp[137]+tmp[38]*tmp[136]+tmp[39]*tmp[135]+tmp[40]*tmp[134]+tmp[41]*tmp[133]+tmp[42]*tmp[132]+tmp[43]*tmp[131]+tmp[44]*tmp[130]+tmp[45]*tmp[129]+tmp[46]*tmp[128]+tmp[47]*tmp[127]+tmp[48]*tmp[126]+tmp[49]*tmp[125]+tmp[50]*tmp[124]+tmp[51]*tmp[123]+tmp[52]*tmp[122]+tmp[53]*tmp[121]+tmp[54]*tmp[120]+tmp[55]*tmp[119]+tmp[56]*tmp[118]+tmp[57]*tmp[117]+tmp[58]*tmp[116]+tmp[59]*tmp[115]+tmp[60]*tmp[114]+tmp[61]*tmp[113]+tmp[62]*tmp[112]+tmp[63]*tmp[111]+tmp[64]*tmp[110]+tmp[65]*tmp[109]+tmp[66]*tmp[108]+tmp[67]*tmp[107]+tmp[68]*tmp[106]+tmp[69]*tmp[105]+tmp[70]*tmp[104]+tmp[71]*tmp[103]+tmp[72]*tmp[102]+tmp[73]*tmp[101]+tmp[74]*tmp[100];
				ans[75]<=tmp[0]*tmp[175]+tmp[1]*tmp[174]+tmp[2]*tmp[173]+tmp[3]*tmp[172]+tmp[4]*tmp[171]+tmp[5]*tmp[170]+tmp[6]*tmp[169]+tmp[7]*tmp[168]+tmp[8]*tmp[167]+tmp[9]*tmp[166]+tmp[10]*tmp[165]+tmp[11]*tmp[164]+tmp[12]*tmp[163]+tmp[13]*tmp[162]+tmp[14]*tmp[161]+tmp[15]*tmp[160]+tmp[16]*tmp[159]+tmp[17]*tmp[158]+tmp[18]*tmp[157]+tmp[19]*tmp[156]+tmp[20]*tmp[155]+tmp[21]*tmp[154]+tmp[22]*tmp[153]+tmp[23]*tmp[152]+tmp[24]*tmp[151]+tmp[25]*tmp[150]+tmp[26]*tmp[149]+tmp[27]*tmp[148]+tmp[28]*tmp[147]+tmp[29]*tmp[146]+tmp[30]*tmp[145]+tmp[31]*tmp[144]+tmp[32]*tmp[143]+tmp[33]*tmp[142]+tmp[34]*tmp[141]+tmp[35]*tmp[140]+tmp[36]*tmp[139]+tmp[37]*tmp[138]+tmp[38]*tmp[137]+tmp[39]*tmp[136]+tmp[40]*tmp[135]+tmp[41]*tmp[134]+tmp[42]*tmp[133]+tmp[43]*tmp[132]+tmp[44]*tmp[131]+tmp[45]*tmp[130]+tmp[46]*tmp[129]+tmp[47]*tmp[128]+tmp[48]*tmp[127]+tmp[49]*tmp[126]+tmp[50]*tmp[125]+tmp[51]*tmp[124]+tmp[52]*tmp[123]+tmp[53]*tmp[122]+tmp[54]*tmp[121]+tmp[55]*tmp[120]+tmp[56]*tmp[119]+tmp[57]*tmp[118]+tmp[58]*tmp[117]+tmp[59]*tmp[116]+tmp[60]*tmp[115]+tmp[61]*tmp[114]+tmp[62]*tmp[113]+tmp[63]*tmp[112]+tmp[64]*tmp[111]+tmp[65]*tmp[110]+tmp[66]*tmp[109]+tmp[67]*tmp[108]+tmp[68]*tmp[107]+tmp[69]*tmp[106]+tmp[70]*tmp[105]+tmp[71]*tmp[104]+tmp[72]*tmp[103]+tmp[73]*tmp[102]+tmp[74]*tmp[101]+tmp[75]*tmp[100];
				ans[76]<=tmp[0]*tmp[176]+tmp[1]*tmp[175]+tmp[2]*tmp[174]+tmp[3]*tmp[173]+tmp[4]*tmp[172]+tmp[5]*tmp[171]+tmp[6]*tmp[170]+tmp[7]*tmp[169]+tmp[8]*tmp[168]+tmp[9]*tmp[167]+tmp[10]*tmp[166]+tmp[11]*tmp[165]+tmp[12]*tmp[164]+tmp[13]*tmp[163]+tmp[14]*tmp[162]+tmp[15]*tmp[161]+tmp[16]*tmp[160]+tmp[17]*tmp[159]+tmp[18]*tmp[158]+tmp[19]*tmp[157]+tmp[20]*tmp[156]+tmp[21]*tmp[155]+tmp[22]*tmp[154]+tmp[23]*tmp[153]+tmp[24]*tmp[152]+tmp[25]*tmp[151]+tmp[26]*tmp[150]+tmp[27]*tmp[149]+tmp[28]*tmp[148]+tmp[29]*tmp[147]+tmp[30]*tmp[146]+tmp[31]*tmp[145]+tmp[32]*tmp[144]+tmp[33]*tmp[143]+tmp[34]*tmp[142]+tmp[35]*tmp[141]+tmp[36]*tmp[140]+tmp[37]*tmp[139]+tmp[38]*tmp[138]+tmp[39]*tmp[137]+tmp[40]*tmp[136]+tmp[41]*tmp[135]+tmp[42]*tmp[134]+tmp[43]*tmp[133]+tmp[44]*tmp[132]+tmp[45]*tmp[131]+tmp[46]*tmp[130]+tmp[47]*tmp[129]+tmp[48]*tmp[128]+tmp[49]*tmp[127]+tmp[50]*tmp[126]+tmp[51]*tmp[125]+tmp[52]*tmp[124]+tmp[53]*tmp[123]+tmp[54]*tmp[122]+tmp[55]*tmp[121]+tmp[56]*tmp[120]+tmp[57]*tmp[119]+tmp[58]*tmp[118]+tmp[59]*tmp[117]+tmp[60]*tmp[116]+tmp[61]*tmp[115]+tmp[62]*tmp[114]+tmp[63]*tmp[113]+tmp[64]*tmp[112]+tmp[65]*tmp[111]+tmp[66]*tmp[110]+tmp[67]*tmp[109]+tmp[68]*tmp[108]+tmp[69]*tmp[107]+tmp[70]*tmp[106]+tmp[71]*tmp[105]+tmp[72]*tmp[104]+tmp[73]*tmp[103]+tmp[74]*tmp[102]+tmp[75]*tmp[101]+tmp[76]*tmp[100];
				ans[77]<=tmp[0]*tmp[177]+tmp[1]*tmp[176]+tmp[2]*tmp[175]+tmp[3]*tmp[174]+tmp[4]*tmp[173]+tmp[5]*tmp[172]+tmp[6]*tmp[171]+tmp[7]*tmp[170]+tmp[8]*tmp[169]+tmp[9]*tmp[168]+tmp[10]*tmp[167]+tmp[11]*tmp[166]+tmp[12]*tmp[165]+tmp[13]*tmp[164]+tmp[14]*tmp[163]+tmp[15]*tmp[162]+tmp[16]*tmp[161]+tmp[17]*tmp[160]+tmp[18]*tmp[159]+tmp[19]*tmp[158]+tmp[20]*tmp[157]+tmp[21]*tmp[156]+tmp[22]*tmp[155]+tmp[23]*tmp[154]+tmp[24]*tmp[153]+tmp[25]*tmp[152]+tmp[26]*tmp[151]+tmp[27]*tmp[150]+tmp[28]*tmp[149]+tmp[29]*tmp[148]+tmp[30]*tmp[147]+tmp[31]*tmp[146]+tmp[32]*tmp[145]+tmp[33]*tmp[144]+tmp[34]*tmp[143]+tmp[35]*tmp[142]+tmp[36]*tmp[141]+tmp[37]*tmp[140]+tmp[38]*tmp[139]+tmp[39]*tmp[138]+tmp[40]*tmp[137]+tmp[41]*tmp[136]+tmp[42]*tmp[135]+tmp[43]*tmp[134]+tmp[44]*tmp[133]+tmp[45]*tmp[132]+tmp[46]*tmp[131]+tmp[47]*tmp[130]+tmp[48]*tmp[129]+tmp[49]*tmp[128]+tmp[50]*tmp[127]+tmp[51]*tmp[126]+tmp[52]*tmp[125]+tmp[53]*tmp[124]+tmp[54]*tmp[123]+tmp[55]*tmp[122]+tmp[56]*tmp[121]+tmp[57]*tmp[120]+tmp[58]*tmp[119]+tmp[59]*tmp[118]+tmp[60]*tmp[117]+tmp[61]*tmp[116]+tmp[62]*tmp[115]+tmp[63]*tmp[114]+tmp[64]*tmp[113]+tmp[65]*tmp[112]+tmp[66]*tmp[111]+tmp[67]*tmp[110]+tmp[68]*tmp[109]+tmp[69]*tmp[108]+tmp[70]*tmp[107]+tmp[71]*tmp[106]+tmp[72]*tmp[105]+tmp[73]*tmp[104]+tmp[74]*tmp[103]+tmp[75]*tmp[102]+tmp[76]*tmp[101]+tmp[77]*tmp[100];
				ans[78]<=tmp[0]*tmp[178]+tmp[1]*tmp[177]+tmp[2]*tmp[176]+tmp[3]*tmp[175]+tmp[4]*tmp[174]+tmp[5]*tmp[173]+tmp[6]*tmp[172]+tmp[7]*tmp[171]+tmp[8]*tmp[170]+tmp[9]*tmp[169]+tmp[10]*tmp[168]+tmp[11]*tmp[167]+tmp[12]*tmp[166]+tmp[13]*tmp[165]+tmp[14]*tmp[164]+tmp[15]*tmp[163]+tmp[16]*tmp[162]+tmp[17]*tmp[161]+tmp[18]*tmp[160]+tmp[19]*tmp[159]+tmp[20]*tmp[158]+tmp[21]*tmp[157]+tmp[22]*tmp[156]+tmp[23]*tmp[155]+tmp[24]*tmp[154]+tmp[25]*tmp[153]+tmp[26]*tmp[152]+tmp[27]*tmp[151]+tmp[28]*tmp[150]+tmp[29]*tmp[149]+tmp[30]*tmp[148]+tmp[31]*tmp[147]+tmp[32]*tmp[146]+tmp[33]*tmp[145]+tmp[34]*tmp[144]+tmp[35]*tmp[143]+tmp[36]*tmp[142]+tmp[37]*tmp[141]+tmp[38]*tmp[140]+tmp[39]*tmp[139]+tmp[40]*tmp[138]+tmp[41]*tmp[137]+tmp[42]*tmp[136]+tmp[43]*tmp[135]+tmp[44]*tmp[134]+tmp[45]*tmp[133]+tmp[46]*tmp[132]+tmp[47]*tmp[131]+tmp[48]*tmp[130]+tmp[49]*tmp[129]+tmp[50]*tmp[128]+tmp[51]*tmp[127]+tmp[52]*tmp[126]+tmp[53]*tmp[125]+tmp[54]*tmp[124]+tmp[55]*tmp[123]+tmp[56]*tmp[122]+tmp[57]*tmp[121]+tmp[58]*tmp[120]+tmp[59]*tmp[119]+tmp[60]*tmp[118]+tmp[61]*tmp[117]+tmp[62]*tmp[116]+tmp[63]*tmp[115]+tmp[64]*tmp[114]+tmp[65]*tmp[113]+tmp[66]*tmp[112]+tmp[67]*tmp[111]+tmp[68]*tmp[110]+tmp[69]*tmp[109]+tmp[70]*tmp[108]+tmp[71]*tmp[107]+tmp[72]*tmp[106]+tmp[73]*tmp[105]+tmp[74]*tmp[104]+tmp[75]*tmp[103]+tmp[76]*tmp[102]+tmp[77]*tmp[101]+tmp[78]*tmp[100];
				ans[79]<=tmp[0]*tmp[179]+tmp[1]*tmp[178]+tmp[2]*tmp[177]+tmp[3]*tmp[176]+tmp[4]*tmp[175]+tmp[5]*tmp[174]+tmp[6]*tmp[173]+tmp[7]*tmp[172]+tmp[8]*tmp[171]+tmp[9]*tmp[170]+tmp[10]*tmp[169]+tmp[11]*tmp[168]+tmp[12]*tmp[167]+tmp[13]*tmp[166]+tmp[14]*tmp[165]+tmp[15]*tmp[164]+tmp[16]*tmp[163]+tmp[17]*tmp[162]+tmp[18]*tmp[161]+tmp[19]*tmp[160]+tmp[20]*tmp[159]+tmp[21]*tmp[158]+tmp[22]*tmp[157]+tmp[23]*tmp[156]+tmp[24]*tmp[155]+tmp[25]*tmp[154]+tmp[26]*tmp[153]+tmp[27]*tmp[152]+tmp[28]*tmp[151]+tmp[29]*tmp[150]+tmp[30]*tmp[149]+tmp[31]*tmp[148]+tmp[32]*tmp[147]+tmp[33]*tmp[146]+tmp[34]*tmp[145]+tmp[35]*tmp[144]+tmp[36]*tmp[143]+tmp[37]*tmp[142]+tmp[38]*tmp[141]+tmp[39]*tmp[140]+tmp[40]*tmp[139]+tmp[41]*tmp[138]+tmp[42]*tmp[137]+tmp[43]*tmp[136]+tmp[44]*tmp[135]+tmp[45]*tmp[134]+tmp[46]*tmp[133]+tmp[47]*tmp[132]+tmp[48]*tmp[131]+tmp[49]*tmp[130]+tmp[50]*tmp[129]+tmp[51]*tmp[128]+tmp[52]*tmp[127]+tmp[53]*tmp[126]+tmp[54]*tmp[125]+tmp[55]*tmp[124]+tmp[56]*tmp[123]+tmp[57]*tmp[122]+tmp[58]*tmp[121]+tmp[59]*tmp[120]+tmp[60]*tmp[119]+tmp[61]*tmp[118]+tmp[62]*tmp[117]+tmp[63]*tmp[116]+tmp[64]*tmp[115]+tmp[65]*tmp[114]+tmp[66]*tmp[113]+tmp[67]*tmp[112]+tmp[68]*tmp[111]+tmp[69]*tmp[110]+tmp[70]*tmp[109]+tmp[71]*tmp[108]+tmp[72]*tmp[107]+tmp[73]*tmp[106]+tmp[74]*tmp[105]+tmp[75]*tmp[104]+tmp[76]*tmp[103]+tmp[77]*tmp[102]+tmp[78]*tmp[101]+tmp[79]*tmp[100];
				ans[80]<=tmp[0]*tmp[180]+tmp[1]*tmp[179]+tmp[2]*tmp[178]+tmp[3]*tmp[177]+tmp[4]*tmp[176]+tmp[5]*tmp[175]+tmp[6]*tmp[174]+tmp[7]*tmp[173]+tmp[8]*tmp[172]+tmp[9]*tmp[171]+tmp[10]*tmp[170]+tmp[11]*tmp[169]+tmp[12]*tmp[168]+tmp[13]*tmp[167]+tmp[14]*tmp[166]+tmp[15]*tmp[165]+tmp[16]*tmp[164]+tmp[17]*tmp[163]+tmp[18]*tmp[162]+tmp[19]*tmp[161]+tmp[20]*tmp[160]+tmp[21]*tmp[159]+tmp[22]*tmp[158]+tmp[23]*tmp[157]+tmp[24]*tmp[156]+tmp[25]*tmp[155]+tmp[26]*tmp[154]+tmp[27]*tmp[153]+tmp[28]*tmp[152]+tmp[29]*tmp[151]+tmp[30]*tmp[150]+tmp[31]*tmp[149]+tmp[32]*tmp[148]+tmp[33]*tmp[147]+tmp[34]*tmp[146]+tmp[35]*tmp[145]+tmp[36]*tmp[144]+tmp[37]*tmp[143]+tmp[38]*tmp[142]+tmp[39]*tmp[141]+tmp[40]*tmp[140]+tmp[41]*tmp[139]+tmp[42]*tmp[138]+tmp[43]*tmp[137]+tmp[44]*tmp[136]+tmp[45]*tmp[135]+tmp[46]*tmp[134]+tmp[47]*tmp[133]+tmp[48]*tmp[132]+tmp[49]*tmp[131]+tmp[50]*tmp[130]+tmp[51]*tmp[129]+tmp[52]*tmp[128]+tmp[53]*tmp[127]+tmp[54]*tmp[126]+tmp[55]*tmp[125]+tmp[56]*tmp[124]+tmp[57]*tmp[123]+tmp[58]*tmp[122]+tmp[59]*tmp[121]+tmp[60]*tmp[120]+tmp[61]*tmp[119]+tmp[62]*tmp[118]+tmp[63]*tmp[117]+tmp[64]*tmp[116]+tmp[65]*tmp[115]+tmp[66]*tmp[114]+tmp[67]*tmp[113]+tmp[68]*tmp[112]+tmp[69]*tmp[111]+tmp[70]*tmp[110]+tmp[71]*tmp[109]+tmp[72]*tmp[108]+tmp[73]*tmp[107]+tmp[74]*tmp[106]+tmp[75]*tmp[105]+tmp[76]*tmp[104]+tmp[77]*tmp[103]+tmp[78]*tmp[102]+tmp[79]*tmp[101]+tmp[80]*tmp[100];
				ans[81]<=tmp[0]*tmp[181]+tmp[1]*tmp[180]+tmp[2]*tmp[179]+tmp[3]*tmp[178]+tmp[4]*tmp[177]+tmp[5]*tmp[176]+tmp[6]*tmp[175]+tmp[7]*tmp[174]+tmp[8]*tmp[173]+tmp[9]*tmp[172]+tmp[10]*tmp[171]+tmp[11]*tmp[170]+tmp[12]*tmp[169]+tmp[13]*tmp[168]+tmp[14]*tmp[167]+tmp[15]*tmp[166]+tmp[16]*tmp[165]+tmp[17]*tmp[164]+tmp[18]*tmp[163]+tmp[19]*tmp[162]+tmp[20]*tmp[161]+tmp[21]*tmp[160]+tmp[22]*tmp[159]+tmp[23]*tmp[158]+tmp[24]*tmp[157]+tmp[25]*tmp[156]+tmp[26]*tmp[155]+tmp[27]*tmp[154]+tmp[28]*tmp[153]+tmp[29]*tmp[152]+tmp[30]*tmp[151]+tmp[31]*tmp[150]+tmp[32]*tmp[149]+tmp[33]*tmp[148]+tmp[34]*tmp[147]+tmp[35]*tmp[146]+tmp[36]*tmp[145]+tmp[37]*tmp[144]+tmp[38]*tmp[143]+tmp[39]*tmp[142]+tmp[40]*tmp[141]+tmp[41]*tmp[140]+tmp[42]*tmp[139]+tmp[43]*tmp[138]+tmp[44]*tmp[137]+tmp[45]*tmp[136]+tmp[46]*tmp[135]+tmp[47]*tmp[134]+tmp[48]*tmp[133]+tmp[49]*tmp[132]+tmp[50]*tmp[131]+tmp[51]*tmp[130]+tmp[52]*tmp[129]+tmp[53]*tmp[128]+tmp[54]*tmp[127]+tmp[55]*tmp[126]+tmp[56]*tmp[125]+tmp[57]*tmp[124]+tmp[58]*tmp[123]+tmp[59]*tmp[122]+tmp[60]*tmp[121]+tmp[61]*tmp[120]+tmp[62]*tmp[119]+tmp[63]*tmp[118]+tmp[64]*tmp[117]+tmp[65]*tmp[116]+tmp[66]*tmp[115]+tmp[67]*tmp[114]+tmp[68]*tmp[113]+tmp[69]*tmp[112]+tmp[70]*tmp[111]+tmp[71]*tmp[110]+tmp[72]*tmp[109]+tmp[73]*tmp[108]+tmp[74]*tmp[107]+tmp[75]*tmp[106]+tmp[76]*tmp[105]+tmp[77]*tmp[104]+tmp[78]*tmp[103]+tmp[79]*tmp[102]+tmp[80]*tmp[101]+tmp[81]*tmp[100];
				ans[82]<=tmp[0]*tmp[182]+tmp[1]*tmp[181]+tmp[2]*tmp[180]+tmp[3]*tmp[179]+tmp[4]*tmp[178]+tmp[5]*tmp[177]+tmp[6]*tmp[176]+tmp[7]*tmp[175]+tmp[8]*tmp[174]+tmp[9]*tmp[173]+tmp[10]*tmp[172]+tmp[11]*tmp[171]+tmp[12]*tmp[170]+tmp[13]*tmp[169]+tmp[14]*tmp[168]+tmp[15]*tmp[167]+tmp[16]*tmp[166]+tmp[17]*tmp[165]+tmp[18]*tmp[164]+tmp[19]*tmp[163]+tmp[20]*tmp[162]+tmp[21]*tmp[161]+tmp[22]*tmp[160]+tmp[23]*tmp[159]+tmp[24]*tmp[158]+tmp[25]*tmp[157]+tmp[26]*tmp[156]+tmp[27]*tmp[155]+tmp[28]*tmp[154]+tmp[29]*tmp[153]+tmp[30]*tmp[152]+tmp[31]*tmp[151]+tmp[32]*tmp[150]+tmp[33]*tmp[149]+tmp[34]*tmp[148]+tmp[35]*tmp[147]+tmp[36]*tmp[146]+tmp[37]*tmp[145]+tmp[38]*tmp[144]+tmp[39]*tmp[143]+tmp[40]*tmp[142]+tmp[41]*tmp[141]+tmp[42]*tmp[140]+tmp[43]*tmp[139]+tmp[44]*tmp[138]+tmp[45]*tmp[137]+tmp[46]*tmp[136]+tmp[47]*tmp[135]+tmp[48]*tmp[134]+tmp[49]*tmp[133]+tmp[50]*tmp[132]+tmp[51]*tmp[131]+tmp[52]*tmp[130]+tmp[53]*tmp[129]+tmp[54]*tmp[128]+tmp[55]*tmp[127]+tmp[56]*tmp[126]+tmp[57]*tmp[125]+tmp[58]*tmp[124]+tmp[59]*tmp[123]+tmp[60]*tmp[122]+tmp[61]*tmp[121]+tmp[62]*tmp[120]+tmp[63]*tmp[119]+tmp[64]*tmp[118]+tmp[65]*tmp[117]+tmp[66]*tmp[116]+tmp[67]*tmp[115]+tmp[68]*tmp[114]+tmp[69]*tmp[113]+tmp[70]*tmp[112]+tmp[71]*tmp[111]+tmp[72]*tmp[110]+tmp[73]*tmp[109]+tmp[74]*tmp[108]+tmp[75]*tmp[107]+tmp[76]*tmp[106]+tmp[77]*tmp[105]+tmp[78]*tmp[104]+tmp[79]*tmp[103]+tmp[80]*tmp[102]+tmp[81]*tmp[101]+tmp[82]*tmp[100];
				ans[83]<=tmp[0]*tmp[183]+tmp[1]*tmp[182]+tmp[2]*tmp[181]+tmp[3]*tmp[180]+tmp[4]*tmp[179]+tmp[5]*tmp[178]+tmp[6]*tmp[177]+tmp[7]*tmp[176]+tmp[8]*tmp[175]+tmp[9]*tmp[174]+tmp[10]*tmp[173]+tmp[11]*tmp[172]+tmp[12]*tmp[171]+tmp[13]*tmp[170]+tmp[14]*tmp[169]+tmp[15]*tmp[168]+tmp[16]*tmp[167]+tmp[17]*tmp[166]+tmp[18]*tmp[165]+tmp[19]*tmp[164]+tmp[20]*tmp[163]+tmp[21]*tmp[162]+tmp[22]*tmp[161]+tmp[23]*tmp[160]+tmp[24]*tmp[159]+tmp[25]*tmp[158]+tmp[26]*tmp[157]+tmp[27]*tmp[156]+tmp[28]*tmp[155]+tmp[29]*tmp[154]+tmp[30]*tmp[153]+tmp[31]*tmp[152]+tmp[32]*tmp[151]+tmp[33]*tmp[150]+tmp[34]*tmp[149]+tmp[35]*tmp[148]+tmp[36]*tmp[147]+tmp[37]*tmp[146]+tmp[38]*tmp[145]+tmp[39]*tmp[144]+tmp[40]*tmp[143]+tmp[41]*tmp[142]+tmp[42]*tmp[141]+tmp[43]*tmp[140]+tmp[44]*tmp[139]+tmp[45]*tmp[138]+tmp[46]*tmp[137]+tmp[47]*tmp[136]+tmp[48]*tmp[135]+tmp[49]*tmp[134]+tmp[50]*tmp[133]+tmp[51]*tmp[132]+tmp[52]*tmp[131]+tmp[53]*tmp[130]+tmp[54]*tmp[129]+tmp[55]*tmp[128]+tmp[56]*tmp[127]+tmp[57]*tmp[126]+tmp[58]*tmp[125]+tmp[59]*tmp[124]+tmp[60]*tmp[123]+tmp[61]*tmp[122]+tmp[62]*tmp[121]+tmp[63]*tmp[120]+tmp[64]*tmp[119]+tmp[65]*tmp[118]+tmp[66]*tmp[117]+tmp[67]*tmp[116]+tmp[68]*tmp[115]+tmp[69]*tmp[114]+tmp[70]*tmp[113]+tmp[71]*tmp[112]+tmp[72]*tmp[111]+tmp[73]*tmp[110]+tmp[74]*tmp[109]+tmp[75]*tmp[108]+tmp[76]*tmp[107]+tmp[77]*tmp[106]+tmp[78]*tmp[105]+tmp[79]*tmp[104]+tmp[80]*tmp[103]+tmp[81]*tmp[102]+tmp[82]*tmp[101]+tmp[83]*tmp[100];
				ans[84]<=tmp[0]*tmp[184]+tmp[1]*tmp[183]+tmp[2]*tmp[182]+tmp[3]*tmp[181]+tmp[4]*tmp[180]+tmp[5]*tmp[179]+tmp[6]*tmp[178]+tmp[7]*tmp[177]+tmp[8]*tmp[176]+tmp[9]*tmp[175]+tmp[10]*tmp[174]+tmp[11]*tmp[173]+tmp[12]*tmp[172]+tmp[13]*tmp[171]+tmp[14]*tmp[170]+tmp[15]*tmp[169]+tmp[16]*tmp[168]+tmp[17]*tmp[167]+tmp[18]*tmp[166]+tmp[19]*tmp[165]+tmp[20]*tmp[164]+tmp[21]*tmp[163]+tmp[22]*tmp[162]+tmp[23]*tmp[161]+tmp[24]*tmp[160]+tmp[25]*tmp[159]+tmp[26]*tmp[158]+tmp[27]*tmp[157]+tmp[28]*tmp[156]+tmp[29]*tmp[155]+tmp[30]*tmp[154]+tmp[31]*tmp[153]+tmp[32]*tmp[152]+tmp[33]*tmp[151]+tmp[34]*tmp[150]+tmp[35]*tmp[149]+tmp[36]*tmp[148]+tmp[37]*tmp[147]+tmp[38]*tmp[146]+tmp[39]*tmp[145]+tmp[40]*tmp[144]+tmp[41]*tmp[143]+tmp[42]*tmp[142]+tmp[43]*tmp[141]+tmp[44]*tmp[140]+tmp[45]*tmp[139]+tmp[46]*tmp[138]+tmp[47]*tmp[137]+tmp[48]*tmp[136]+tmp[49]*tmp[135]+tmp[50]*tmp[134]+tmp[51]*tmp[133]+tmp[52]*tmp[132]+tmp[53]*tmp[131]+tmp[54]*tmp[130]+tmp[55]*tmp[129]+tmp[56]*tmp[128]+tmp[57]*tmp[127]+tmp[58]*tmp[126]+tmp[59]*tmp[125]+tmp[60]*tmp[124]+tmp[61]*tmp[123]+tmp[62]*tmp[122]+tmp[63]*tmp[121]+tmp[64]*tmp[120]+tmp[65]*tmp[119]+tmp[66]*tmp[118]+tmp[67]*tmp[117]+tmp[68]*tmp[116]+tmp[69]*tmp[115]+tmp[70]*tmp[114]+tmp[71]*tmp[113]+tmp[72]*tmp[112]+tmp[73]*tmp[111]+tmp[74]*tmp[110]+tmp[75]*tmp[109]+tmp[76]*tmp[108]+tmp[77]*tmp[107]+tmp[78]*tmp[106]+tmp[79]*tmp[105]+tmp[80]*tmp[104]+tmp[81]*tmp[103]+tmp[82]*tmp[102]+tmp[83]*tmp[101]+tmp[84]*tmp[100];
				ans[85]<=tmp[0]*tmp[185]+tmp[1]*tmp[184]+tmp[2]*tmp[183]+tmp[3]*tmp[182]+tmp[4]*tmp[181]+tmp[5]*tmp[180]+tmp[6]*tmp[179]+tmp[7]*tmp[178]+tmp[8]*tmp[177]+tmp[9]*tmp[176]+tmp[10]*tmp[175]+tmp[11]*tmp[174]+tmp[12]*tmp[173]+tmp[13]*tmp[172]+tmp[14]*tmp[171]+tmp[15]*tmp[170]+tmp[16]*tmp[169]+tmp[17]*tmp[168]+tmp[18]*tmp[167]+tmp[19]*tmp[166]+tmp[20]*tmp[165]+tmp[21]*tmp[164]+tmp[22]*tmp[163]+tmp[23]*tmp[162]+tmp[24]*tmp[161]+tmp[25]*tmp[160]+tmp[26]*tmp[159]+tmp[27]*tmp[158]+tmp[28]*tmp[157]+tmp[29]*tmp[156]+tmp[30]*tmp[155]+tmp[31]*tmp[154]+tmp[32]*tmp[153]+tmp[33]*tmp[152]+tmp[34]*tmp[151]+tmp[35]*tmp[150]+tmp[36]*tmp[149]+tmp[37]*tmp[148]+tmp[38]*tmp[147]+tmp[39]*tmp[146]+tmp[40]*tmp[145]+tmp[41]*tmp[144]+tmp[42]*tmp[143]+tmp[43]*tmp[142]+tmp[44]*tmp[141]+tmp[45]*tmp[140]+tmp[46]*tmp[139]+tmp[47]*tmp[138]+tmp[48]*tmp[137]+tmp[49]*tmp[136]+tmp[50]*tmp[135]+tmp[51]*tmp[134]+tmp[52]*tmp[133]+tmp[53]*tmp[132]+tmp[54]*tmp[131]+tmp[55]*tmp[130]+tmp[56]*tmp[129]+tmp[57]*tmp[128]+tmp[58]*tmp[127]+tmp[59]*tmp[126]+tmp[60]*tmp[125]+tmp[61]*tmp[124]+tmp[62]*tmp[123]+tmp[63]*tmp[122]+tmp[64]*tmp[121]+tmp[65]*tmp[120]+tmp[66]*tmp[119]+tmp[67]*tmp[118]+tmp[68]*tmp[117]+tmp[69]*tmp[116]+tmp[70]*tmp[115]+tmp[71]*tmp[114]+tmp[72]*tmp[113]+tmp[73]*tmp[112]+tmp[74]*tmp[111]+tmp[75]*tmp[110]+tmp[76]*tmp[109]+tmp[77]*tmp[108]+tmp[78]*tmp[107]+tmp[79]*tmp[106]+tmp[80]*tmp[105]+tmp[81]*tmp[104]+tmp[82]*tmp[103]+tmp[83]*tmp[102]+tmp[84]*tmp[101]+tmp[85]*tmp[100];
				ans[86]<=tmp[0]*tmp[186]+tmp[1]*tmp[185]+tmp[2]*tmp[184]+tmp[3]*tmp[183]+tmp[4]*tmp[182]+tmp[5]*tmp[181]+tmp[6]*tmp[180]+tmp[7]*tmp[179]+tmp[8]*tmp[178]+tmp[9]*tmp[177]+tmp[10]*tmp[176]+tmp[11]*tmp[175]+tmp[12]*tmp[174]+tmp[13]*tmp[173]+tmp[14]*tmp[172]+tmp[15]*tmp[171]+tmp[16]*tmp[170]+tmp[17]*tmp[169]+tmp[18]*tmp[168]+tmp[19]*tmp[167]+tmp[20]*tmp[166]+tmp[21]*tmp[165]+tmp[22]*tmp[164]+tmp[23]*tmp[163]+tmp[24]*tmp[162]+tmp[25]*tmp[161]+tmp[26]*tmp[160]+tmp[27]*tmp[159]+tmp[28]*tmp[158]+tmp[29]*tmp[157]+tmp[30]*tmp[156]+tmp[31]*tmp[155]+tmp[32]*tmp[154]+tmp[33]*tmp[153]+tmp[34]*tmp[152]+tmp[35]*tmp[151]+tmp[36]*tmp[150]+tmp[37]*tmp[149]+tmp[38]*tmp[148]+tmp[39]*tmp[147]+tmp[40]*tmp[146]+tmp[41]*tmp[145]+tmp[42]*tmp[144]+tmp[43]*tmp[143]+tmp[44]*tmp[142]+tmp[45]*tmp[141]+tmp[46]*tmp[140]+tmp[47]*tmp[139]+tmp[48]*tmp[138]+tmp[49]*tmp[137]+tmp[50]*tmp[136]+tmp[51]*tmp[135]+tmp[52]*tmp[134]+tmp[53]*tmp[133]+tmp[54]*tmp[132]+tmp[55]*tmp[131]+tmp[56]*tmp[130]+tmp[57]*tmp[129]+tmp[58]*tmp[128]+tmp[59]*tmp[127]+tmp[60]*tmp[126]+tmp[61]*tmp[125]+tmp[62]*tmp[124]+tmp[63]*tmp[123]+tmp[64]*tmp[122]+tmp[65]*tmp[121]+tmp[66]*tmp[120]+tmp[67]*tmp[119]+tmp[68]*tmp[118]+tmp[69]*tmp[117]+tmp[70]*tmp[116]+tmp[71]*tmp[115]+tmp[72]*tmp[114]+tmp[73]*tmp[113]+tmp[74]*tmp[112]+tmp[75]*tmp[111]+tmp[76]*tmp[110]+tmp[77]*tmp[109]+tmp[78]*tmp[108]+tmp[79]*tmp[107]+tmp[80]*tmp[106]+tmp[81]*tmp[105]+tmp[82]*tmp[104]+tmp[83]*tmp[103]+tmp[84]*tmp[102]+tmp[85]*tmp[101]+tmp[86]*tmp[100];
				ans[87]<=tmp[0]*tmp[187]+tmp[1]*tmp[186]+tmp[2]*tmp[185]+tmp[3]*tmp[184]+tmp[4]*tmp[183]+tmp[5]*tmp[182]+tmp[6]*tmp[181]+tmp[7]*tmp[180]+tmp[8]*tmp[179]+tmp[9]*tmp[178]+tmp[10]*tmp[177]+tmp[11]*tmp[176]+tmp[12]*tmp[175]+tmp[13]*tmp[174]+tmp[14]*tmp[173]+tmp[15]*tmp[172]+tmp[16]*tmp[171]+tmp[17]*tmp[170]+tmp[18]*tmp[169]+tmp[19]*tmp[168]+tmp[20]*tmp[167]+tmp[21]*tmp[166]+tmp[22]*tmp[165]+tmp[23]*tmp[164]+tmp[24]*tmp[163]+tmp[25]*tmp[162]+tmp[26]*tmp[161]+tmp[27]*tmp[160]+tmp[28]*tmp[159]+tmp[29]*tmp[158]+tmp[30]*tmp[157]+tmp[31]*tmp[156]+tmp[32]*tmp[155]+tmp[33]*tmp[154]+tmp[34]*tmp[153]+tmp[35]*tmp[152]+tmp[36]*tmp[151]+tmp[37]*tmp[150]+tmp[38]*tmp[149]+tmp[39]*tmp[148]+tmp[40]*tmp[147]+tmp[41]*tmp[146]+tmp[42]*tmp[145]+tmp[43]*tmp[144]+tmp[44]*tmp[143]+tmp[45]*tmp[142]+tmp[46]*tmp[141]+tmp[47]*tmp[140]+tmp[48]*tmp[139]+tmp[49]*tmp[138]+tmp[50]*tmp[137]+tmp[51]*tmp[136]+tmp[52]*tmp[135]+tmp[53]*tmp[134]+tmp[54]*tmp[133]+tmp[55]*tmp[132]+tmp[56]*tmp[131]+tmp[57]*tmp[130]+tmp[58]*tmp[129]+tmp[59]*tmp[128]+tmp[60]*tmp[127]+tmp[61]*tmp[126]+tmp[62]*tmp[125]+tmp[63]*tmp[124]+tmp[64]*tmp[123]+tmp[65]*tmp[122]+tmp[66]*tmp[121]+tmp[67]*tmp[120]+tmp[68]*tmp[119]+tmp[69]*tmp[118]+tmp[70]*tmp[117]+tmp[71]*tmp[116]+tmp[72]*tmp[115]+tmp[73]*tmp[114]+tmp[74]*tmp[113]+tmp[75]*tmp[112]+tmp[76]*tmp[111]+tmp[77]*tmp[110]+tmp[78]*tmp[109]+tmp[79]*tmp[108]+tmp[80]*tmp[107]+tmp[81]*tmp[106]+tmp[82]*tmp[105]+tmp[83]*tmp[104]+tmp[84]*tmp[103]+tmp[85]*tmp[102]+tmp[86]*tmp[101]+tmp[87]*tmp[100];
				ans[88]<=tmp[0]*tmp[188]+tmp[1]*tmp[187]+tmp[2]*tmp[186]+tmp[3]*tmp[185]+tmp[4]*tmp[184]+tmp[5]*tmp[183]+tmp[6]*tmp[182]+tmp[7]*tmp[181]+tmp[8]*tmp[180]+tmp[9]*tmp[179]+tmp[10]*tmp[178]+tmp[11]*tmp[177]+tmp[12]*tmp[176]+tmp[13]*tmp[175]+tmp[14]*tmp[174]+tmp[15]*tmp[173]+tmp[16]*tmp[172]+tmp[17]*tmp[171]+tmp[18]*tmp[170]+tmp[19]*tmp[169]+tmp[20]*tmp[168]+tmp[21]*tmp[167]+tmp[22]*tmp[166]+tmp[23]*tmp[165]+tmp[24]*tmp[164]+tmp[25]*tmp[163]+tmp[26]*tmp[162]+tmp[27]*tmp[161]+tmp[28]*tmp[160]+tmp[29]*tmp[159]+tmp[30]*tmp[158]+tmp[31]*tmp[157]+tmp[32]*tmp[156]+tmp[33]*tmp[155]+tmp[34]*tmp[154]+tmp[35]*tmp[153]+tmp[36]*tmp[152]+tmp[37]*tmp[151]+tmp[38]*tmp[150]+tmp[39]*tmp[149]+tmp[40]*tmp[148]+tmp[41]*tmp[147]+tmp[42]*tmp[146]+tmp[43]*tmp[145]+tmp[44]*tmp[144]+tmp[45]*tmp[143]+tmp[46]*tmp[142]+tmp[47]*tmp[141]+tmp[48]*tmp[140]+tmp[49]*tmp[139]+tmp[50]*tmp[138]+tmp[51]*tmp[137]+tmp[52]*tmp[136]+tmp[53]*tmp[135]+tmp[54]*tmp[134]+tmp[55]*tmp[133]+tmp[56]*tmp[132]+tmp[57]*tmp[131]+tmp[58]*tmp[130]+tmp[59]*tmp[129]+tmp[60]*tmp[128]+tmp[61]*tmp[127]+tmp[62]*tmp[126]+tmp[63]*tmp[125]+tmp[64]*tmp[124]+tmp[65]*tmp[123]+tmp[66]*tmp[122]+tmp[67]*tmp[121]+tmp[68]*tmp[120]+tmp[69]*tmp[119]+tmp[70]*tmp[118]+tmp[71]*tmp[117]+tmp[72]*tmp[116]+tmp[73]*tmp[115]+tmp[74]*tmp[114]+tmp[75]*tmp[113]+tmp[76]*tmp[112]+tmp[77]*tmp[111]+tmp[78]*tmp[110]+tmp[79]*tmp[109]+tmp[80]*tmp[108]+tmp[81]*tmp[107]+tmp[82]*tmp[106]+tmp[83]*tmp[105]+tmp[84]*tmp[104]+tmp[85]*tmp[103]+tmp[86]*tmp[102]+tmp[87]*tmp[101]+tmp[88]*tmp[100];
				ans[89]<=tmp[0]*tmp[189]+tmp[1]*tmp[188]+tmp[2]*tmp[187]+tmp[3]*tmp[186]+tmp[4]*tmp[185]+tmp[5]*tmp[184]+tmp[6]*tmp[183]+tmp[7]*tmp[182]+tmp[8]*tmp[181]+tmp[9]*tmp[180]+tmp[10]*tmp[179]+tmp[11]*tmp[178]+tmp[12]*tmp[177]+tmp[13]*tmp[176]+tmp[14]*tmp[175]+tmp[15]*tmp[174]+tmp[16]*tmp[173]+tmp[17]*tmp[172]+tmp[18]*tmp[171]+tmp[19]*tmp[170]+tmp[20]*tmp[169]+tmp[21]*tmp[168]+tmp[22]*tmp[167]+tmp[23]*tmp[166]+tmp[24]*tmp[165]+tmp[25]*tmp[164]+tmp[26]*tmp[163]+tmp[27]*tmp[162]+tmp[28]*tmp[161]+tmp[29]*tmp[160]+tmp[30]*tmp[159]+tmp[31]*tmp[158]+tmp[32]*tmp[157]+tmp[33]*tmp[156]+tmp[34]*tmp[155]+tmp[35]*tmp[154]+tmp[36]*tmp[153]+tmp[37]*tmp[152]+tmp[38]*tmp[151]+tmp[39]*tmp[150]+tmp[40]*tmp[149]+tmp[41]*tmp[148]+tmp[42]*tmp[147]+tmp[43]*tmp[146]+tmp[44]*tmp[145]+tmp[45]*tmp[144]+tmp[46]*tmp[143]+tmp[47]*tmp[142]+tmp[48]*tmp[141]+tmp[49]*tmp[140]+tmp[50]*tmp[139]+tmp[51]*tmp[138]+tmp[52]*tmp[137]+tmp[53]*tmp[136]+tmp[54]*tmp[135]+tmp[55]*tmp[134]+tmp[56]*tmp[133]+tmp[57]*tmp[132]+tmp[58]*tmp[131]+tmp[59]*tmp[130]+tmp[60]*tmp[129]+tmp[61]*tmp[128]+tmp[62]*tmp[127]+tmp[63]*tmp[126]+tmp[64]*tmp[125]+tmp[65]*tmp[124]+tmp[66]*tmp[123]+tmp[67]*tmp[122]+tmp[68]*tmp[121]+tmp[69]*tmp[120]+tmp[70]*tmp[119]+tmp[71]*tmp[118]+tmp[72]*tmp[117]+tmp[73]*tmp[116]+tmp[74]*tmp[115]+tmp[75]*tmp[114]+tmp[76]*tmp[113]+tmp[77]*tmp[112]+tmp[78]*tmp[111]+tmp[79]*tmp[110]+tmp[80]*tmp[109]+tmp[81]*tmp[108]+tmp[82]*tmp[107]+tmp[83]*tmp[106]+tmp[84]*tmp[105]+tmp[85]*tmp[104]+tmp[86]*tmp[103]+tmp[87]*tmp[102]+tmp[88]*tmp[101]+tmp[89]*tmp[100];
				ans[90]<=tmp[0]*tmp[190]+tmp[1]*tmp[189]+tmp[2]*tmp[188]+tmp[3]*tmp[187]+tmp[4]*tmp[186]+tmp[5]*tmp[185]+tmp[6]*tmp[184]+tmp[7]*tmp[183]+tmp[8]*tmp[182]+tmp[9]*tmp[181]+tmp[10]*tmp[180]+tmp[11]*tmp[179]+tmp[12]*tmp[178]+tmp[13]*tmp[177]+tmp[14]*tmp[176]+tmp[15]*tmp[175]+tmp[16]*tmp[174]+tmp[17]*tmp[173]+tmp[18]*tmp[172]+tmp[19]*tmp[171]+tmp[20]*tmp[170]+tmp[21]*tmp[169]+tmp[22]*tmp[168]+tmp[23]*tmp[167]+tmp[24]*tmp[166]+tmp[25]*tmp[165]+tmp[26]*tmp[164]+tmp[27]*tmp[163]+tmp[28]*tmp[162]+tmp[29]*tmp[161]+tmp[30]*tmp[160]+tmp[31]*tmp[159]+tmp[32]*tmp[158]+tmp[33]*tmp[157]+tmp[34]*tmp[156]+tmp[35]*tmp[155]+tmp[36]*tmp[154]+tmp[37]*tmp[153]+tmp[38]*tmp[152]+tmp[39]*tmp[151]+tmp[40]*tmp[150]+tmp[41]*tmp[149]+tmp[42]*tmp[148]+tmp[43]*tmp[147]+tmp[44]*tmp[146]+tmp[45]*tmp[145]+tmp[46]*tmp[144]+tmp[47]*tmp[143]+tmp[48]*tmp[142]+tmp[49]*tmp[141]+tmp[50]*tmp[140]+tmp[51]*tmp[139]+tmp[52]*tmp[138]+tmp[53]*tmp[137]+tmp[54]*tmp[136]+tmp[55]*tmp[135]+tmp[56]*tmp[134]+tmp[57]*tmp[133]+tmp[58]*tmp[132]+tmp[59]*tmp[131]+tmp[60]*tmp[130]+tmp[61]*tmp[129]+tmp[62]*tmp[128]+tmp[63]*tmp[127]+tmp[64]*tmp[126]+tmp[65]*tmp[125]+tmp[66]*tmp[124]+tmp[67]*tmp[123]+tmp[68]*tmp[122]+tmp[69]*tmp[121]+tmp[70]*tmp[120]+tmp[71]*tmp[119]+tmp[72]*tmp[118]+tmp[73]*tmp[117]+tmp[74]*tmp[116]+tmp[75]*tmp[115]+tmp[76]*tmp[114]+tmp[77]*tmp[113]+tmp[78]*tmp[112]+tmp[79]*tmp[111]+tmp[80]*tmp[110]+tmp[81]*tmp[109]+tmp[82]*tmp[108]+tmp[83]*tmp[107]+tmp[84]*tmp[106]+tmp[85]*tmp[105]+tmp[86]*tmp[104]+tmp[87]*tmp[103]+tmp[88]*tmp[102]+tmp[89]*tmp[101]+tmp[90]*tmp[100];
				ans[91]<=tmp[0]*tmp[191]+tmp[1]*tmp[190]+tmp[2]*tmp[189]+tmp[3]*tmp[188]+tmp[4]*tmp[187]+tmp[5]*tmp[186]+tmp[6]*tmp[185]+tmp[7]*tmp[184]+tmp[8]*tmp[183]+tmp[9]*tmp[182]+tmp[10]*tmp[181]+tmp[11]*tmp[180]+tmp[12]*tmp[179]+tmp[13]*tmp[178]+tmp[14]*tmp[177]+tmp[15]*tmp[176]+tmp[16]*tmp[175]+tmp[17]*tmp[174]+tmp[18]*tmp[173]+tmp[19]*tmp[172]+tmp[20]*tmp[171]+tmp[21]*tmp[170]+tmp[22]*tmp[169]+tmp[23]*tmp[168]+tmp[24]*tmp[167]+tmp[25]*tmp[166]+tmp[26]*tmp[165]+tmp[27]*tmp[164]+tmp[28]*tmp[163]+tmp[29]*tmp[162]+tmp[30]*tmp[161]+tmp[31]*tmp[160]+tmp[32]*tmp[159]+tmp[33]*tmp[158]+tmp[34]*tmp[157]+tmp[35]*tmp[156]+tmp[36]*tmp[155]+tmp[37]*tmp[154]+tmp[38]*tmp[153]+tmp[39]*tmp[152]+tmp[40]*tmp[151]+tmp[41]*tmp[150]+tmp[42]*tmp[149]+tmp[43]*tmp[148]+tmp[44]*tmp[147]+tmp[45]*tmp[146]+tmp[46]*tmp[145]+tmp[47]*tmp[144]+tmp[48]*tmp[143]+tmp[49]*tmp[142]+tmp[50]*tmp[141]+tmp[51]*tmp[140]+tmp[52]*tmp[139]+tmp[53]*tmp[138]+tmp[54]*tmp[137]+tmp[55]*tmp[136]+tmp[56]*tmp[135]+tmp[57]*tmp[134]+tmp[58]*tmp[133]+tmp[59]*tmp[132]+tmp[60]*tmp[131]+tmp[61]*tmp[130]+tmp[62]*tmp[129]+tmp[63]*tmp[128]+tmp[64]*tmp[127]+tmp[65]*tmp[126]+tmp[66]*tmp[125]+tmp[67]*tmp[124]+tmp[68]*tmp[123]+tmp[69]*tmp[122]+tmp[70]*tmp[121]+tmp[71]*tmp[120]+tmp[72]*tmp[119]+tmp[73]*tmp[118]+tmp[74]*tmp[117]+tmp[75]*tmp[116]+tmp[76]*tmp[115]+tmp[77]*tmp[114]+tmp[78]*tmp[113]+tmp[79]*tmp[112]+tmp[80]*tmp[111]+tmp[81]*tmp[110]+tmp[82]*tmp[109]+tmp[83]*tmp[108]+tmp[84]*tmp[107]+tmp[85]*tmp[106]+tmp[86]*tmp[105]+tmp[87]*tmp[104]+tmp[88]*tmp[103]+tmp[89]*tmp[102]+tmp[90]*tmp[101]+tmp[91]*tmp[100];
				ans[92]<=tmp[0]*tmp[192]+tmp[1]*tmp[191]+tmp[2]*tmp[190]+tmp[3]*tmp[189]+tmp[4]*tmp[188]+tmp[5]*tmp[187]+tmp[6]*tmp[186]+tmp[7]*tmp[185]+tmp[8]*tmp[184]+tmp[9]*tmp[183]+tmp[10]*tmp[182]+tmp[11]*tmp[181]+tmp[12]*tmp[180]+tmp[13]*tmp[179]+tmp[14]*tmp[178]+tmp[15]*tmp[177]+tmp[16]*tmp[176]+tmp[17]*tmp[175]+tmp[18]*tmp[174]+tmp[19]*tmp[173]+tmp[20]*tmp[172]+tmp[21]*tmp[171]+tmp[22]*tmp[170]+tmp[23]*tmp[169]+tmp[24]*tmp[168]+tmp[25]*tmp[167]+tmp[26]*tmp[166]+tmp[27]*tmp[165]+tmp[28]*tmp[164]+tmp[29]*tmp[163]+tmp[30]*tmp[162]+tmp[31]*tmp[161]+tmp[32]*tmp[160]+tmp[33]*tmp[159]+tmp[34]*tmp[158]+tmp[35]*tmp[157]+tmp[36]*tmp[156]+tmp[37]*tmp[155]+tmp[38]*tmp[154]+tmp[39]*tmp[153]+tmp[40]*tmp[152]+tmp[41]*tmp[151]+tmp[42]*tmp[150]+tmp[43]*tmp[149]+tmp[44]*tmp[148]+tmp[45]*tmp[147]+tmp[46]*tmp[146]+tmp[47]*tmp[145]+tmp[48]*tmp[144]+tmp[49]*tmp[143]+tmp[50]*tmp[142]+tmp[51]*tmp[141]+tmp[52]*tmp[140]+tmp[53]*tmp[139]+tmp[54]*tmp[138]+tmp[55]*tmp[137]+tmp[56]*tmp[136]+tmp[57]*tmp[135]+tmp[58]*tmp[134]+tmp[59]*tmp[133]+tmp[60]*tmp[132]+tmp[61]*tmp[131]+tmp[62]*tmp[130]+tmp[63]*tmp[129]+tmp[64]*tmp[128]+tmp[65]*tmp[127]+tmp[66]*tmp[126]+tmp[67]*tmp[125]+tmp[68]*tmp[124]+tmp[69]*tmp[123]+tmp[70]*tmp[122]+tmp[71]*tmp[121]+tmp[72]*tmp[120]+tmp[73]*tmp[119]+tmp[74]*tmp[118]+tmp[75]*tmp[117]+tmp[76]*tmp[116]+tmp[77]*tmp[115]+tmp[78]*tmp[114]+tmp[79]*tmp[113]+tmp[80]*tmp[112]+tmp[81]*tmp[111]+tmp[82]*tmp[110]+tmp[83]*tmp[109]+tmp[84]*tmp[108]+tmp[85]*tmp[107]+tmp[86]*tmp[106]+tmp[87]*tmp[105]+tmp[88]*tmp[104]+tmp[89]*tmp[103]+tmp[90]*tmp[102]+tmp[91]*tmp[101]+tmp[92]*tmp[100];
				ans[93]<=tmp[0]*tmp[193]+tmp[1]*tmp[192]+tmp[2]*tmp[191]+tmp[3]*tmp[190]+tmp[4]*tmp[189]+tmp[5]*tmp[188]+tmp[6]*tmp[187]+tmp[7]*tmp[186]+tmp[8]*tmp[185]+tmp[9]*tmp[184]+tmp[10]*tmp[183]+tmp[11]*tmp[182]+tmp[12]*tmp[181]+tmp[13]*tmp[180]+tmp[14]*tmp[179]+tmp[15]*tmp[178]+tmp[16]*tmp[177]+tmp[17]*tmp[176]+tmp[18]*tmp[175]+tmp[19]*tmp[174]+tmp[20]*tmp[173]+tmp[21]*tmp[172]+tmp[22]*tmp[171]+tmp[23]*tmp[170]+tmp[24]*tmp[169]+tmp[25]*tmp[168]+tmp[26]*tmp[167]+tmp[27]*tmp[166]+tmp[28]*tmp[165]+tmp[29]*tmp[164]+tmp[30]*tmp[163]+tmp[31]*tmp[162]+tmp[32]*tmp[161]+tmp[33]*tmp[160]+tmp[34]*tmp[159]+tmp[35]*tmp[158]+tmp[36]*tmp[157]+tmp[37]*tmp[156]+tmp[38]*tmp[155]+tmp[39]*tmp[154]+tmp[40]*tmp[153]+tmp[41]*tmp[152]+tmp[42]*tmp[151]+tmp[43]*tmp[150]+tmp[44]*tmp[149]+tmp[45]*tmp[148]+tmp[46]*tmp[147]+tmp[47]*tmp[146]+tmp[48]*tmp[145]+tmp[49]*tmp[144]+tmp[50]*tmp[143]+tmp[51]*tmp[142]+tmp[52]*tmp[141]+tmp[53]*tmp[140]+tmp[54]*tmp[139]+tmp[55]*tmp[138]+tmp[56]*tmp[137]+tmp[57]*tmp[136]+tmp[58]*tmp[135]+tmp[59]*tmp[134]+tmp[60]*tmp[133]+tmp[61]*tmp[132]+tmp[62]*tmp[131]+tmp[63]*tmp[130]+tmp[64]*tmp[129]+tmp[65]*tmp[128]+tmp[66]*tmp[127]+tmp[67]*tmp[126]+tmp[68]*tmp[125]+tmp[69]*tmp[124]+tmp[70]*tmp[123]+tmp[71]*tmp[122]+tmp[72]*tmp[121]+tmp[73]*tmp[120]+tmp[74]*tmp[119]+tmp[75]*tmp[118]+tmp[76]*tmp[117]+tmp[77]*tmp[116]+tmp[78]*tmp[115]+tmp[79]*tmp[114]+tmp[80]*tmp[113]+tmp[81]*tmp[112]+tmp[82]*tmp[111]+tmp[83]*tmp[110]+tmp[84]*tmp[109]+tmp[85]*tmp[108]+tmp[86]*tmp[107]+tmp[87]*tmp[106]+tmp[88]*tmp[105]+tmp[89]*tmp[104]+tmp[90]*tmp[103]+tmp[91]*tmp[102]+tmp[92]*tmp[101]+tmp[93]*tmp[100];
				ans[94]<=tmp[0]*tmp[194]+tmp[1]*tmp[193]+tmp[2]*tmp[192]+tmp[3]*tmp[191]+tmp[4]*tmp[190]+tmp[5]*tmp[189]+tmp[6]*tmp[188]+tmp[7]*tmp[187]+tmp[8]*tmp[186]+tmp[9]*tmp[185]+tmp[10]*tmp[184]+tmp[11]*tmp[183]+tmp[12]*tmp[182]+tmp[13]*tmp[181]+tmp[14]*tmp[180]+tmp[15]*tmp[179]+tmp[16]*tmp[178]+tmp[17]*tmp[177]+tmp[18]*tmp[176]+tmp[19]*tmp[175]+tmp[20]*tmp[174]+tmp[21]*tmp[173]+tmp[22]*tmp[172]+tmp[23]*tmp[171]+tmp[24]*tmp[170]+tmp[25]*tmp[169]+tmp[26]*tmp[168]+tmp[27]*tmp[167]+tmp[28]*tmp[166]+tmp[29]*tmp[165]+tmp[30]*tmp[164]+tmp[31]*tmp[163]+tmp[32]*tmp[162]+tmp[33]*tmp[161]+tmp[34]*tmp[160]+tmp[35]*tmp[159]+tmp[36]*tmp[158]+tmp[37]*tmp[157]+tmp[38]*tmp[156]+tmp[39]*tmp[155]+tmp[40]*tmp[154]+tmp[41]*tmp[153]+tmp[42]*tmp[152]+tmp[43]*tmp[151]+tmp[44]*tmp[150]+tmp[45]*tmp[149]+tmp[46]*tmp[148]+tmp[47]*tmp[147]+tmp[48]*tmp[146]+tmp[49]*tmp[145]+tmp[50]*tmp[144]+tmp[51]*tmp[143]+tmp[52]*tmp[142]+tmp[53]*tmp[141]+tmp[54]*tmp[140]+tmp[55]*tmp[139]+tmp[56]*tmp[138]+tmp[57]*tmp[137]+tmp[58]*tmp[136]+tmp[59]*tmp[135]+tmp[60]*tmp[134]+tmp[61]*tmp[133]+tmp[62]*tmp[132]+tmp[63]*tmp[131]+tmp[64]*tmp[130]+tmp[65]*tmp[129]+tmp[66]*tmp[128]+tmp[67]*tmp[127]+tmp[68]*tmp[126]+tmp[69]*tmp[125]+tmp[70]*tmp[124]+tmp[71]*tmp[123]+tmp[72]*tmp[122]+tmp[73]*tmp[121]+tmp[74]*tmp[120]+tmp[75]*tmp[119]+tmp[76]*tmp[118]+tmp[77]*tmp[117]+tmp[78]*tmp[116]+tmp[79]*tmp[115]+tmp[80]*tmp[114]+tmp[81]*tmp[113]+tmp[82]*tmp[112]+tmp[83]*tmp[111]+tmp[84]*tmp[110]+tmp[85]*tmp[109]+tmp[86]*tmp[108]+tmp[87]*tmp[107]+tmp[88]*tmp[106]+tmp[89]*tmp[105]+tmp[90]*tmp[104]+tmp[91]*tmp[103]+tmp[92]*tmp[102]+tmp[93]*tmp[101]+tmp[94]*tmp[100];
				ans[95]<=tmp[0]*tmp[195]+tmp[1]*tmp[194]+tmp[2]*tmp[193]+tmp[3]*tmp[192]+tmp[4]*tmp[191]+tmp[5]*tmp[190]+tmp[6]*tmp[189]+tmp[7]*tmp[188]+tmp[8]*tmp[187]+tmp[9]*tmp[186]+tmp[10]*tmp[185]+tmp[11]*tmp[184]+tmp[12]*tmp[183]+tmp[13]*tmp[182]+tmp[14]*tmp[181]+tmp[15]*tmp[180]+tmp[16]*tmp[179]+tmp[17]*tmp[178]+tmp[18]*tmp[177]+tmp[19]*tmp[176]+tmp[20]*tmp[175]+tmp[21]*tmp[174]+tmp[22]*tmp[173]+tmp[23]*tmp[172]+tmp[24]*tmp[171]+tmp[25]*tmp[170]+tmp[26]*tmp[169]+tmp[27]*tmp[168]+tmp[28]*tmp[167]+tmp[29]*tmp[166]+tmp[30]*tmp[165]+tmp[31]*tmp[164]+tmp[32]*tmp[163]+tmp[33]*tmp[162]+tmp[34]*tmp[161]+tmp[35]*tmp[160]+tmp[36]*tmp[159]+tmp[37]*tmp[158]+tmp[38]*tmp[157]+tmp[39]*tmp[156]+tmp[40]*tmp[155]+tmp[41]*tmp[154]+tmp[42]*tmp[153]+tmp[43]*tmp[152]+tmp[44]*tmp[151]+tmp[45]*tmp[150]+tmp[46]*tmp[149]+tmp[47]*tmp[148]+tmp[48]*tmp[147]+tmp[49]*tmp[146]+tmp[50]*tmp[145]+tmp[51]*tmp[144]+tmp[52]*tmp[143]+tmp[53]*tmp[142]+tmp[54]*tmp[141]+tmp[55]*tmp[140]+tmp[56]*tmp[139]+tmp[57]*tmp[138]+tmp[58]*tmp[137]+tmp[59]*tmp[136]+tmp[60]*tmp[135]+tmp[61]*tmp[134]+tmp[62]*tmp[133]+tmp[63]*tmp[132]+tmp[64]*tmp[131]+tmp[65]*tmp[130]+tmp[66]*tmp[129]+tmp[67]*tmp[128]+tmp[68]*tmp[127]+tmp[69]*tmp[126]+tmp[70]*tmp[125]+tmp[71]*tmp[124]+tmp[72]*tmp[123]+tmp[73]*tmp[122]+tmp[74]*tmp[121]+tmp[75]*tmp[120]+tmp[76]*tmp[119]+tmp[77]*tmp[118]+tmp[78]*tmp[117]+tmp[79]*tmp[116]+tmp[80]*tmp[115]+tmp[81]*tmp[114]+tmp[82]*tmp[113]+tmp[83]*tmp[112]+tmp[84]*tmp[111]+tmp[85]*tmp[110]+tmp[86]*tmp[109]+tmp[87]*tmp[108]+tmp[88]*tmp[107]+tmp[89]*tmp[106]+tmp[90]*tmp[105]+tmp[91]*tmp[104]+tmp[92]*tmp[103]+tmp[93]*tmp[102]+tmp[94]*tmp[101]+tmp[95]*tmp[100];
				ans[96]<=tmp[0]*tmp[196]+tmp[1]*tmp[195]+tmp[2]*tmp[194]+tmp[3]*tmp[193]+tmp[4]*tmp[192]+tmp[5]*tmp[191]+tmp[6]*tmp[190]+tmp[7]*tmp[189]+tmp[8]*tmp[188]+tmp[9]*tmp[187]+tmp[10]*tmp[186]+tmp[11]*tmp[185]+tmp[12]*tmp[184]+tmp[13]*tmp[183]+tmp[14]*tmp[182]+tmp[15]*tmp[181]+tmp[16]*tmp[180]+tmp[17]*tmp[179]+tmp[18]*tmp[178]+tmp[19]*tmp[177]+tmp[20]*tmp[176]+tmp[21]*tmp[175]+tmp[22]*tmp[174]+tmp[23]*tmp[173]+tmp[24]*tmp[172]+tmp[25]*tmp[171]+tmp[26]*tmp[170]+tmp[27]*tmp[169]+tmp[28]*tmp[168]+tmp[29]*tmp[167]+tmp[30]*tmp[166]+tmp[31]*tmp[165]+tmp[32]*tmp[164]+tmp[33]*tmp[163]+tmp[34]*tmp[162]+tmp[35]*tmp[161]+tmp[36]*tmp[160]+tmp[37]*tmp[159]+tmp[38]*tmp[158]+tmp[39]*tmp[157]+tmp[40]*tmp[156]+tmp[41]*tmp[155]+tmp[42]*tmp[154]+tmp[43]*tmp[153]+tmp[44]*tmp[152]+tmp[45]*tmp[151]+tmp[46]*tmp[150]+tmp[47]*tmp[149]+tmp[48]*tmp[148]+tmp[49]*tmp[147]+tmp[50]*tmp[146]+tmp[51]*tmp[145]+tmp[52]*tmp[144]+tmp[53]*tmp[143]+tmp[54]*tmp[142]+tmp[55]*tmp[141]+tmp[56]*tmp[140]+tmp[57]*tmp[139]+tmp[58]*tmp[138]+tmp[59]*tmp[137]+tmp[60]*tmp[136]+tmp[61]*tmp[135]+tmp[62]*tmp[134]+tmp[63]*tmp[133]+tmp[64]*tmp[132]+tmp[65]*tmp[131]+tmp[66]*tmp[130]+tmp[67]*tmp[129]+tmp[68]*tmp[128]+tmp[69]*tmp[127]+tmp[70]*tmp[126]+tmp[71]*tmp[125]+tmp[72]*tmp[124]+tmp[73]*tmp[123]+tmp[74]*tmp[122]+tmp[75]*tmp[121]+tmp[76]*tmp[120]+tmp[77]*tmp[119]+tmp[78]*tmp[118]+tmp[79]*tmp[117]+tmp[80]*tmp[116]+tmp[81]*tmp[115]+tmp[82]*tmp[114]+tmp[83]*tmp[113]+tmp[84]*tmp[112]+tmp[85]*tmp[111]+tmp[86]*tmp[110]+tmp[87]*tmp[109]+tmp[88]*tmp[108]+tmp[89]*tmp[107]+tmp[90]*tmp[106]+tmp[91]*tmp[105]+tmp[92]*tmp[104]+tmp[93]*tmp[103]+tmp[94]*tmp[102]+tmp[95]*tmp[101]+tmp[96]*tmp[100];
				ans[97]<=tmp[0]*tmp[197]+tmp[1]*tmp[196]+tmp[2]*tmp[195]+tmp[3]*tmp[194]+tmp[4]*tmp[193]+tmp[5]*tmp[192]+tmp[6]*tmp[191]+tmp[7]*tmp[190]+tmp[8]*tmp[189]+tmp[9]*tmp[188]+tmp[10]*tmp[187]+tmp[11]*tmp[186]+tmp[12]*tmp[185]+tmp[13]*tmp[184]+tmp[14]*tmp[183]+tmp[15]*tmp[182]+tmp[16]*tmp[181]+tmp[17]*tmp[180]+tmp[18]*tmp[179]+tmp[19]*tmp[178]+tmp[20]*tmp[177]+tmp[21]*tmp[176]+tmp[22]*tmp[175]+tmp[23]*tmp[174]+tmp[24]*tmp[173]+tmp[25]*tmp[172]+tmp[26]*tmp[171]+tmp[27]*tmp[170]+tmp[28]*tmp[169]+tmp[29]*tmp[168]+tmp[30]*tmp[167]+tmp[31]*tmp[166]+tmp[32]*tmp[165]+tmp[33]*tmp[164]+tmp[34]*tmp[163]+tmp[35]*tmp[162]+tmp[36]*tmp[161]+tmp[37]*tmp[160]+tmp[38]*tmp[159]+tmp[39]*tmp[158]+tmp[40]*tmp[157]+tmp[41]*tmp[156]+tmp[42]*tmp[155]+tmp[43]*tmp[154]+tmp[44]*tmp[153]+tmp[45]*tmp[152]+tmp[46]*tmp[151]+tmp[47]*tmp[150]+tmp[48]*tmp[149]+tmp[49]*tmp[148]+tmp[50]*tmp[147]+tmp[51]*tmp[146]+tmp[52]*tmp[145]+tmp[53]*tmp[144]+tmp[54]*tmp[143]+tmp[55]*tmp[142]+tmp[56]*tmp[141]+tmp[57]*tmp[140]+tmp[58]*tmp[139]+tmp[59]*tmp[138]+tmp[60]*tmp[137]+tmp[61]*tmp[136]+tmp[62]*tmp[135]+tmp[63]*tmp[134]+tmp[64]*tmp[133]+tmp[65]*tmp[132]+tmp[66]*tmp[131]+tmp[67]*tmp[130]+tmp[68]*tmp[129]+tmp[69]*tmp[128]+tmp[70]*tmp[127]+tmp[71]*tmp[126]+tmp[72]*tmp[125]+tmp[73]*tmp[124]+tmp[74]*tmp[123]+tmp[75]*tmp[122]+tmp[76]*tmp[121]+tmp[77]*tmp[120]+tmp[78]*tmp[119]+tmp[79]*tmp[118]+tmp[80]*tmp[117]+tmp[81]*tmp[116]+tmp[82]*tmp[115]+tmp[83]*tmp[114]+tmp[84]*tmp[113]+tmp[85]*tmp[112]+tmp[86]*tmp[111]+tmp[87]*tmp[110]+tmp[88]*tmp[109]+tmp[89]*tmp[108]+tmp[90]*tmp[107]+tmp[91]*tmp[106]+tmp[92]*tmp[105]+tmp[93]*tmp[104]+tmp[94]*tmp[103]+tmp[95]*tmp[102]+tmp[96]*tmp[101]+tmp[97]*tmp[100];
				ans[98]<=tmp[0]*tmp[198]+tmp[1]*tmp[197]+tmp[2]*tmp[196]+tmp[3]*tmp[195]+tmp[4]*tmp[194]+tmp[5]*tmp[193]+tmp[6]*tmp[192]+tmp[7]*tmp[191]+tmp[8]*tmp[190]+tmp[9]*tmp[189]+tmp[10]*tmp[188]+tmp[11]*tmp[187]+tmp[12]*tmp[186]+tmp[13]*tmp[185]+tmp[14]*tmp[184]+tmp[15]*tmp[183]+tmp[16]*tmp[182]+tmp[17]*tmp[181]+tmp[18]*tmp[180]+tmp[19]*tmp[179]+tmp[20]*tmp[178]+tmp[21]*tmp[177]+tmp[22]*tmp[176]+tmp[23]*tmp[175]+tmp[24]*tmp[174]+tmp[25]*tmp[173]+tmp[26]*tmp[172]+tmp[27]*tmp[171]+tmp[28]*tmp[170]+tmp[29]*tmp[169]+tmp[30]*tmp[168]+tmp[31]*tmp[167]+tmp[32]*tmp[166]+tmp[33]*tmp[165]+tmp[34]*tmp[164]+tmp[35]*tmp[163]+tmp[36]*tmp[162]+tmp[37]*tmp[161]+tmp[38]*tmp[160]+tmp[39]*tmp[159]+tmp[40]*tmp[158]+tmp[41]*tmp[157]+tmp[42]*tmp[156]+tmp[43]*tmp[155]+tmp[44]*tmp[154]+tmp[45]*tmp[153]+tmp[46]*tmp[152]+tmp[47]*tmp[151]+tmp[48]*tmp[150]+tmp[49]*tmp[149]+tmp[50]*tmp[148]+tmp[51]*tmp[147]+tmp[52]*tmp[146]+tmp[53]*tmp[145]+tmp[54]*tmp[144]+tmp[55]*tmp[143]+tmp[56]*tmp[142]+tmp[57]*tmp[141]+tmp[58]*tmp[140]+tmp[59]*tmp[139]+tmp[60]*tmp[138]+tmp[61]*tmp[137]+tmp[62]*tmp[136]+tmp[63]*tmp[135]+tmp[64]*tmp[134]+tmp[65]*tmp[133]+tmp[66]*tmp[132]+tmp[67]*tmp[131]+tmp[68]*tmp[130]+tmp[69]*tmp[129]+tmp[70]*tmp[128]+tmp[71]*tmp[127]+tmp[72]*tmp[126]+tmp[73]*tmp[125]+tmp[74]*tmp[124]+tmp[75]*tmp[123]+tmp[76]*tmp[122]+tmp[77]*tmp[121]+tmp[78]*tmp[120]+tmp[79]*tmp[119]+tmp[80]*tmp[118]+tmp[81]*tmp[117]+tmp[82]*tmp[116]+tmp[83]*tmp[115]+tmp[84]*tmp[114]+tmp[85]*tmp[113]+tmp[86]*tmp[112]+tmp[87]*tmp[111]+tmp[88]*tmp[110]+tmp[89]*tmp[109]+tmp[90]*tmp[108]+tmp[91]*tmp[107]+tmp[92]*tmp[106]+tmp[93]*tmp[105]+tmp[94]*tmp[104]+tmp[95]*tmp[103]+tmp[96]*tmp[102]+tmp[97]*tmp[101]+tmp[98]*tmp[100];
				ans[99]<=tmp[0]*tmp[199]+tmp[1]*tmp[198]+tmp[2]*tmp[197]+tmp[3]*tmp[196]+tmp[4]*tmp[195]+tmp[5]*tmp[194]+tmp[6]*tmp[193]+tmp[7]*tmp[192]+tmp[8]*tmp[191]+tmp[9]*tmp[190]+tmp[10]*tmp[189]+tmp[11]*tmp[188]+tmp[12]*tmp[187]+tmp[13]*tmp[186]+tmp[14]*tmp[185]+tmp[15]*tmp[184]+tmp[16]*tmp[183]+tmp[17]*tmp[182]+tmp[18]*tmp[181]+tmp[19]*tmp[180]+tmp[20]*tmp[179]+tmp[21]*tmp[178]+tmp[22]*tmp[177]+tmp[23]*tmp[176]+tmp[24]*tmp[175]+tmp[25]*tmp[174]+tmp[26]*tmp[173]+tmp[27]*tmp[172]+tmp[28]*tmp[171]+tmp[29]*tmp[170]+tmp[30]*tmp[169]+tmp[31]*tmp[168]+tmp[32]*tmp[167]+tmp[33]*tmp[166]+tmp[34]*tmp[165]+tmp[35]*tmp[164]+tmp[36]*tmp[163]+tmp[37]*tmp[162]+tmp[38]*tmp[161]+tmp[39]*tmp[160]+tmp[40]*tmp[159]+tmp[41]*tmp[158]+tmp[42]*tmp[157]+tmp[43]*tmp[156]+tmp[44]*tmp[155]+tmp[45]*tmp[154]+tmp[46]*tmp[153]+tmp[47]*tmp[152]+tmp[48]*tmp[151]+tmp[49]*tmp[150]+tmp[50]*tmp[149]+tmp[51]*tmp[148]+tmp[52]*tmp[147]+tmp[53]*tmp[146]+tmp[54]*tmp[145]+tmp[55]*tmp[144]+tmp[56]*tmp[143]+tmp[57]*tmp[142]+tmp[58]*tmp[141]+tmp[59]*tmp[140]+tmp[60]*tmp[139]+tmp[61]*tmp[138]+tmp[62]*tmp[137]+tmp[63]*tmp[136]+tmp[64]*tmp[135]+tmp[65]*tmp[134]+tmp[66]*tmp[133]+tmp[67]*tmp[132]+tmp[68]*tmp[131]+tmp[69]*tmp[130]+tmp[70]*tmp[129]+tmp[71]*tmp[128]+tmp[72]*tmp[127]+tmp[73]*tmp[126]+tmp[74]*tmp[125]+tmp[75]*tmp[124]+tmp[76]*tmp[123]+tmp[77]*tmp[122]+tmp[78]*tmp[121]+tmp[79]*tmp[120]+tmp[80]*tmp[119]+tmp[81]*tmp[118]+tmp[82]*tmp[117]+tmp[83]*tmp[116]+tmp[84]*tmp[115]+tmp[85]*tmp[114]+tmp[86]*tmp[113]+tmp[87]*tmp[112]+tmp[88]*tmp[111]+tmp[89]*tmp[110]+tmp[90]*tmp[109]+tmp[91]*tmp[108]+tmp[92]*tmp[107]+tmp[93]*tmp[106]+tmp[94]*tmp[105]+tmp[95]*tmp[104]+tmp[96]*tmp[103]+tmp[97]*tmp[102]+tmp[98]*tmp[101]+tmp[99]*tmp[100];
				ans[100]<=tmp[1]*tmp[199]+tmp[2]*tmp[198]+tmp[3]*tmp[197]+tmp[4]*tmp[196]+tmp[5]*tmp[195]+tmp[6]*tmp[194]+tmp[7]*tmp[193]+tmp[8]*tmp[192]+tmp[9]*tmp[191]+tmp[10]*tmp[190]+tmp[11]*tmp[189]+tmp[12]*tmp[188]+tmp[13]*tmp[187]+tmp[14]*tmp[186]+tmp[15]*tmp[185]+tmp[16]*tmp[184]+tmp[17]*tmp[183]+tmp[18]*tmp[182]+tmp[19]*tmp[181]+tmp[20]*tmp[180]+tmp[21]*tmp[179]+tmp[22]*tmp[178]+tmp[23]*tmp[177]+tmp[24]*tmp[176]+tmp[25]*tmp[175]+tmp[26]*tmp[174]+tmp[27]*tmp[173]+tmp[28]*tmp[172]+tmp[29]*tmp[171]+tmp[30]*tmp[170]+tmp[31]*tmp[169]+tmp[32]*tmp[168]+tmp[33]*tmp[167]+tmp[34]*tmp[166]+tmp[35]*tmp[165]+tmp[36]*tmp[164]+tmp[37]*tmp[163]+tmp[38]*tmp[162]+tmp[39]*tmp[161]+tmp[40]*tmp[160]+tmp[41]*tmp[159]+tmp[42]*tmp[158]+tmp[43]*tmp[157]+tmp[44]*tmp[156]+tmp[45]*tmp[155]+tmp[46]*tmp[154]+tmp[47]*tmp[153]+tmp[48]*tmp[152]+tmp[49]*tmp[151]+tmp[50]*tmp[150]+tmp[51]*tmp[149]+tmp[52]*tmp[148]+tmp[53]*tmp[147]+tmp[54]*tmp[146]+tmp[55]*tmp[145]+tmp[56]*tmp[144]+tmp[57]*tmp[143]+tmp[58]*tmp[142]+tmp[59]*tmp[141]+tmp[60]*tmp[140]+tmp[61]*tmp[139]+tmp[62]*tmp[138]+tmp[63]*tmp[137]+tmp[64]*tmp[136]+tmp[65]*tmp[135]+tmp[66]*tmp[134]+tmp[67]*tmp[133]+tmp[68]*tmp[132]+tmp[69]*tmp[131]+tmp[70]*tmp[130]+tmp[71]*tmp[129]+tmp[72]*tmp[128]+tmp[73]*tmp[127]+tmp[74]*tmp[126]+tmp[75]*tmp[125]+tmp[76]*tmp[124]+tmp[77]*tmp[123]+tmp[78]*tmp[122]+tmp[79]*tmp[121]+tmp[80]*tmp[120]+tmp[81]*tmp[119]+tmp[82]*tmp[118]+tmp[83]*tmp[117]+tmp[84]*tmp[116]+tmp[85]*tmp[115]+tmp[86]*tmp[114]+tmp[87]*tmp[113]+tmp[88]*tmp[112]+tmp[89]*tmp[111]+tmp[90]*tmp[110]+tmp[91]*tmp[109]+tmp[92]*tmp[108]+tmp[93]*tmp[107]+tmp[94]*tmp[106]+tmp[95]*tmp[105]+tmp[96]*tmp[104]+tmp[97]*tmp[103]+tmp[98]*tmp[102]+tmp[99]*tmp[101];
				ans[101]<=tmp[2]*tmp[199]+tmp[3]*tmp[198]+tmp[4]*tmp[197]+tmp[5]*tmp[196]+tmp[6]*tmp[195]+tmp[7]*tmp[194]+tmp[8]*tmp[193]+tmp[9]*tmp[192]+tmp[10]*tmp[191]+tmp[11]*tmp[190]+tmp[12]*tmp[189]+tmp[13]*tmp[188]+tmp[14]*tmp[187]+tmp[15]*tmp[186]+tmp[16]*tmp[185]+tmp[17]*tmp[184]+tmp[18]*tmp[183]+tmp[19]*tmp[182]+tmp[20]*tmp[181]+tmp[21]*tmp[180]+tmp[22]*tmp[179]+tmp[23]*tmp[178]+tmp[24]*tmp[177]+tmp[25]*tmp[176]+tmp[26]*tmp[175]+tmp[27]*tmp[174]+tmp[28]*tmp[173]+tmp[29]*tmp[172]+tmp[30]*tmp[171]+tmp[31]*tmp[170]+tmp[32]*tmp[169]+tmp[33]*tmp[168]+tmp[34]*tmp[167]+tmp[35]*tmp[166]+tmp[36]*tmp[165]+tmp[37]*tmp[164]+tmp[38]*tmp[163]+tmp[39]*tmp[162]+tmp[40]*tmp[161]+tmp[41]*tmp[160]+tmp[42]*tmp[159]+tmp[43]*tmp[158]+tmp[44]*tmp[157]+tmp[45]*tmp[156]+tmp[46]*tmp[155]+tmp[47]*tmp[154]+tmp[48]*tmp[153]+tmp[49]*tmp[152]+tmp[50]*tmp[151]+tmp[51]*tmp[150]+tmp[52]*tmp[149]+tmp[53]*tmp[148]+tmp[54]*tmp[147]+tmp[55]*tmp[146]+tmp[56]*tmp[145]+tmp[57]*tmp[144]+tmp[58]*tmp[143]+tmp[59]*tmp[142]+tmp[60]*tmp[141]+tmp[61]*tmp[140]+tmp[62]*tmp[139]+tmp[63]*tmp[138]+tmp[64]*tmp[137]+tmp[65]*tmp[136]+tmp[66]*tmp[135]+tmp[67]*tmp[134]+tmp[68]*tmp[133]+tmp[69]*tmp[132]+tmp[70]*tmp[131]+tmp[71]*tmp[130]+tmp[72]*tmp[129]+tmp[73]*tmp[128]+tmp[74]*tmp[127]+tmp[75]*tmp[126]+tmp[76]*tmp[125]+tmp[77]*tmp[124]+tmp[78]*tmp[123]+tmp[79]*tmp[122]+tmp[80]*tmp[121]+tmp[81]*tmp[120]+tmp[82]*tmp[119]+tmp[83]*tmp[118]+tmp[84]*tmp[117]+tmp[85]*tmp[116]+tmp[86]*tmp[115]+tmp[87]*tmp[114]+tmp[88]*tmp[113]+tmp[89]*tmp[112]+tmp[90]*tmp[111]+tmp[91]*tmp[110]+tmp[92]*tmp[109]+tmp[93]*tmp[108]+tmp[94]*tmp[107]+tmp[95]*tmp[106]+tmp[96]*tmp[105]+tmp[97]*tmp[104]+tmp[98]*tmp[103]+tmp[99]*tmp[102];
				ans[102]<=tmp[3]*tmp[199]+tmp[4]*tmp[198]+tmp[5]*tmp[197]+tmp[6]*tmp[196]+tmp[7]*tmp[195]+tmp[8]*tmp[194]+tmp[9]*tmp[193]+tmp[10]*tmp[192]+tmp[11]*tmp[191]+tmp[12]*tmp[190]+tmp[13]*tmp[189]+tmp[14]*tmp[188]+tmp[15]*tmp[187]+tmp[16]*tmp[186]+tmp[17]*tmp[185]+tmp[18]*tmp[184]+tmp[19]*tmp[183]+tmp[20]*tmp[182]+tmp[21]*tmp[181]+tmp[22]*tmp[180]+tmp[23]*tmp[179]+tmp[24]*tmp[178]+tmp[25]*tmp[177]+tmp[26]*tmp[176]+tmp[27]*tmp[175]+tmp[28]*tmp[174]+tmp[29]*tmp[173]+tmp[30]*tmp[172]+tmp[31]*tmp[171]+tmp[32]*tmp[170]+tmp[33]*tmp[169]+tmp[34]*tmp[168]+tmp[35]*tmp[167]+tmp[36]*tmp[166]+tmp[37]*tmp[165]+tmp[38]*tmp[164]+tmp[39]*tmp[163]+tmp[40]*tmp[162]+tmp[41]*tmp[161]+tmp[42]*tmp[160]+tmp[43]*tmp[159]+tmp[44]*tmp[158]+tmp[45]*tmp[157]+tmp[46]*tmp[156]+tmp[47]*tmp[155]+tmp[48]*tmp[154]+tmp[49]*tmp[153]+tmp[50]*tmp[152]+tmp[51]*tmp[151]+tmp[52]*tmp[150]+tmp[53]*tmp[149]+tmp[54]*tmp[148]+tmp[55]*tmp[147]+tmp[56]*tmp[146]+tmp[57]*tmp[145]+tmp[58]*tmp[144]+tmp[59]*tmp[143]+tmp[60]*tmp[142]+tmp[61]*tmp[141]+tmp[62]*tmp[140]+tmp[63]*tmp[139]+tmp[64]*tmp[138]+tmp[65]*tmp[137]+tmp[66]*tmp[136]+tmp[67]*tmp[135]+tmp[68]*tmp[134]+tmp[69]*tmp[133]+tmp[70]*tmp[132]+tmp[71]*tmp[131]+tmp[72]*tmp[130]+tmp[73]*tmp[129]+tmp[74]*tmp[128]+tmp[75]*tmp[127]+tmp[76]*tmp[126]+tmp[77]*tmp[125]+tmp[78]*tmp[124]+tmp[79]*tmp[123]+tmp[80]*tmp[122]+tmp[81]*tmp[121]+tmp[82]*tmp[120]+tmp[83]*tmp[119]+tmp[84]*tmp[118]+tmp[85]*tmp[117]+tmp[86]*tmp[116]+tmp[87]*tmp[115]+tmp[88]*tmp[114]+tmp[89]*tmp[113]+tmp[90]*tmp[112]+tmp[91]*tmp[111]+tmp[92]*tmp[110]+tmp[93]*tmp[109]+tmp[94]*tmp[108]+tmp[95]*tmp[107]+tmp[96]*tmp[106]+tmp[97]*tmp[105]+tmp[98]*tmp[104]+tmp[99]*tmp[103];
				ans[103]<=tmp[4]*tmp[199]+tmp[5]*tmp[198]+tmp[6]*tmp[197]+tmp[7]*tmp[196]+tmp[8]*tmp[195]+tmp[9]*tmp[194]+tmp[10]*tmp[193]+tmp[11]*tmp[192]+tmp[12]*tmp[191]+tmp[13]*tmp[190]+tmp[14]*tmp[189]+tmp[15]*tmp[188]+tmp[16]*tmp[187]+tmp[17]*tmp[186]+tmp[18]*tmp[185]+tmp[19]*tmp[184]+tmp[20]*tmp[183]+tmp[21]*tmp[182]+tmp[22]*tmp[181]+tmp[23]*tmp[180]+tmp[24]*tmp[179]+tmp[25]*tmp[178]+tmp[26]*tmp[177]+tmp[27]*tmp[176]+tmp[28]*tmp[175]+tmp[29]*tmp[174]+tmp[30]*tmp[173]+tmp[31]*tmp[172]+tmp[32]*tmp[171]+tmp[33]*tmp[170]+tmp[34]*tmp[169]+tmp[35]*tmp[168]+tmp[36]*tmp[167]+tmp[37]*tmp[166]+tmp[38]*tmp[165]+tmp[39]*tmp[164]+tmp[40]*tmp[163]+tmp[41]*tmp[162]+tmp[42]*tmp[161]+tmp[43]*tmp[160]+tmp[44]*tmp[159]+tmp[45]*tmp[158]+tmp[46]*tmp[157]+tmp[47]*tmp[156]+tmp[48]*tmp[155]+tmp[49]*tmp[154]+tmp[50]*tmp[153]+tmp[51]*tmp[152]+tmp[52]*tmp[151]+tmp[53]*tmp[150]+tmp[54]*tmp[149]+tmp[55]*tmp[148]+tmp[56]*tmp[147]+tmp[57]*tmp[146]+tmp[58]*tmp[145]+tmp[59]*tmp[144]+tmp[60]*tmp[143]+tmp[61]*tmp[142]+tmp[62]*tmp[141]+tmp[63]*tmp[140]+tmp[64]*tmp[139]+tmp[65]*tmp[138]+tmp[66]*tmp[137]+tmp[67]*tmp[136]+tmp[68]*tmp[135]+tmp[69]*tmp[134]+tmp[70]*tmp[133]+tmp[71]*tmp[132]+tmp[72]*tmp[131]+tmp[73]*tmp[130]+tmp[74]*tmp[129]+tmp[75]*tmp[128]+tmp[76]*tmp[127]+tmp[77]*tmp[126]+tmp[78]*tmp[125]+tmp[79]*tmp[124]+tmp[80]*tmp[123]+tmp[81]*tmp[122]+tmp[82]*tmp[121]+tmp[83]*tmp[120]+tmp[84]*tmp[119]+tmp[85]*tmp[118]+tmp[86]*tmp[117]+tmp[87]*tmp[116]+tmp[88]*tmp[115]+tmp[89]*tmp[114]+tmp[90]*tmp[113]+tmp[91]*tmp[112]+tmp[92]*tmp[111]+tmp[93]*tmp[110]+tmp[94]*tmp[109]+tmp[95]*tmp[108]+tmp[96]*tmp[107]+tmp[97]*tmp[106]+tmp[98]*tmp[105]+tmp[99]*tmp[104];
				ans[104]<=tmp[5]*tmp[199]+tmp[6]*tmp[198]+tmp[7]*tmp[197]+tmp[8]*tmp[196]+tmp[9]*tmp[195]+tmp[10]*tmp[194]+tmp[11]*tmp[193]+tmp[12]*tmp[192]+tmp[13]*tmp[191]+tmp[14]*tmp[190]+tmp[15]*tmp[189]+tmp[16]*tmp[188]+tmp[17]*tmp[187]+tmp[18]*tmp[186]+tmp[19]*tmp[185]+tmp[20]*tmp[184]+tmp[21]*tmp[183]+tmp[22]*tmp[182]+tmp[23]*tmp[181]+tmp[24]*tmp[180]+tmp[25]*tmp[179]+tmp[26]*tmp[178]+tmp[27]*tmp[177]+tmp[28]*tmp[176]+tmp[29]*tmp[175]+tmp[30]*tmp[174]+tmp[31]*tmp[173]+tmp[32]*tmp[172]+tmp[33]*tmp[171]+tmp[34]*tmp[170]+tmp[35]*tmp[169]+tmp[36]*tmp[168]+tmp[37]*tmp[167]+tmp[38]*tmp[166]+tmp[39]*tmp[165]+tmp[40]*tmp[164]+tmp[41]*tmp[163]+tmp[42]*tmp[162]+tmp[43]*tmp[161]+tmp[44]*tmp[160]+tmp[45]*tmp[159]+tmp[46]*tmp[158]+tmp[47]*tmp[157]+tmp[48]*tmp[156]+tmp[49]*tmp[155]+tmp[50]*tmp[154]+tmp[51]*tmp[153]+tmp[52]*tmp[152]+tmp[53]*tmp[151]+tmp[54]*tmp[150]+tmp[55]*tmp[149]+tmp[56]*tmp[148]+tmp[57]*tmp[147]+tmp[58]*tmp[146]+tmp[59]*tmp[145]+tmp[60]*tmp[144]+tmp[61]*tmp[143]+tmp[62]*tmp[142]+tmp[63]*tmp[141]+tmp[64]*tmp[140]+tmp[65]*tmp[139]+tmp[66]*tmp[138]+tmp[67]*tmp[137]+tmp[68]*tmp[136]+tmp[69]*tmp[135]+tmp[70]*tmp[134]+tmp[71]*tmp[133]+tmp[72]*tmp[132]+tmp[73]*tmp[131]+tmp[74]*tmp[130]+tmp[75]*tmp[129]+tmp[76]*tmp[128]+tmp[77]*tmp[127]+tmp[78]*tmp[126]+tmp[79]*tmp[125]+tmp[80]*tmp[124]+tmp[81]*tmp[123]+tmp[82]*tmp[122]+tmp[83]*tmp[121]+tmp[84]*tmp[120]+tmp[85]*tmp[119]+tmp[86]*tmp[118]+tmp[87]*tmp[117]+tmp[88]*tmp[116]+tmp[89]*tmp[115]+tmp[90]*tmp[114]+tmp[91]*tmp[113]+tmp[92]*tmp[112]+tmp[93]*tmp[111]+tmp[94]*tmp[110]+tmp[95]*tmp[109]+tmp[96]*tmp[108]+tmp[97]*tmp[107]+tmp[98]*tmp[106]+tmp[99]*tmp[105];
				ans[105]<=tmp[6]*tmp[199]+tmp[7]*tmp[198]+tmp[8]*tmp[197]+tmp[9]*tmp[196]+tmp[10]*tmp[195]+tmp[11]*tmp[194]+tmp[12]*tmp[193]+tmp[13]*tmp[192]+tmp[14]*tmp[191]+tmp[15]*tmp[190]+tmp[16]*tmp[189]+tmp[17]*tmp[188]+tmp[18]*tmp[187]+tmp[19]*tmp[186]+tmp[20]*tmp[185]+tmp[21]*tmp[184]+tmp[22]*tmp[183]+tmp[23]*tmp[182]+tmp[24]*tmp[181]+tmp[25]*tmp[180]+tmp[26]*tmp[179]+tmp[27]*tmp[178]+tmp[28]*tmp[177]+tmp[29]*tmp[176]+tmp[30]*tmp[175]+tmp[31]*tmp[174]+tmp[32]*tmp[173]+tmp[33]*tmp[172]+tmp[34]*tmp[171]+tmp[35]*tmp[170]+tmp[36]*tmp[169]+tmp[37]*tmp[168]+tmp[38]*tmp[167]+tmp[39]*tmp[166]+tmp[40]*tmp[165]+tmp[41]*tmp[164]+tmp[42]*tmp[163]+tmp[43]*tmp[162]+tmp[44]*tmp[161]+tmp[45]*tmp[160]+tmp[46]*tmp[159]+tmp[47]*tmp[158]+tmp[48]*tmp[157]+tmp[49]*tmp[156]+tmp[50]*tmp[155]+tmp[51]*tmp[154]+tmp[52]*tmp[153]+tmp[53]*tmp[152]+tmp[54]*tmp[151]+tmp[55]*tmp[150]+tmp[56]*tmp[149]+tmp[57]*tmp[148]+tmp[58]*tmp[147]+tmp[59]*tmp[146]+tmp[60]*tmp[145]+tmp[61]*tmp[144]+tmp[62]*tmp[143]+tmp[63]*tmp[142]+tmp[64]*tmp[141]+tmp[65]*tmp[140]+tmp[66]*tmp[139]+tmp[67]*tmp[138]+tmp[68]*tmp[137]+tmp[69]*tmp[136]+tmp[70]*tmp[135]+tmp[71]*tmp[134]+tmp[72]*tmp[133]+tmp[73]*tmp[132]+tmp[74]*tmp[131]+tmp[75]*tmp[130]+tmp[76]*tmp[129]+tmp[77]*tmp[128]+tmp[78]*tmp[127]+tmp[79]*tmp[126]+tmp[80]*tmp[125]+tmp[81]*tmp[124]+tmp[82]*tmp[123]+tmp[83]*tmp[122]+tmp[84]*tmp[121]+tmp[85]*tmp[120]+tmp[86]*tmp[119]+tmp[87]*tmp[118]+tmp[88]*tmp[117]+tmp[89]*tmp[116]+tmp[90]*tmp[115]+tmp[91]*tmp[114]+tmp[92]*tmp[113]+tmp[93]*tmp[112]+tmp[94]*tmp[111]+tmp[95]*tmp[110]+tmp[96]*tmp[109]+tmp[97]*tmp[108]+tmp[98]*tmp[107]+tmp[99]*tmp[106];
				ans[106]<=tmp[7]*tmp[199]+tmp[8]*tmp[198]+tmp[9]*tmp[197]+tmp[10]*tmp[196]+tmp[11]*tmp[195]+tmp[12]*tmp[194]+tmp[13]*tmp[193]+tmp[14]*tmp[192]+tmp[15]*tmp[191]+tmp[16]*tmp[190]+tmp[17]*tmp[189]+tmp[18]*tmp[188]+tmp[19]*tmp[187]+tmp[20]*tmp[186]+tmp[21]*tmp[185]+tmp[22]*tmp[184]+tmp[23]*tmp[183]+tmp[24]*tmp[182]+tmp[25]*tmp[181]+tmp[26]*tmp[180]+tmp[27]*tmp[179]+tmp[28]*tmp[178]+tmp[29]*tmp[177]+tmp[30]*tmp[176]+tmp[31]*tmp[175]+tmp[32]*tmp[174]+tmp[33]*tmp[173]+tmp[34]*tmp[172]+tmp[35]*tmp[171]+tmp[36]*tmp[170]+tmp[37]*tmp[169]+tmp[38]*tmp[168]+tmp[39]*tmp[167]+tmp[40]*tmp[166]+tmp[41]*tmp[165]+tmp[42]*tmp[164]+tmp[43]*tmp[163]+tmp[44]*tmp[162]+tmp[45]*tmp[161]+tmp[46]*tmp[160]+tmp[47]*tmp[159]+tmp[48]*tmp[158]+tmp[49]*tmp[157]+tmp[50]*tmp[156]+tmp[51]*tmp[155]+tmp[52]*tmp[154]+tmp[53]*tmp[153]+tmp[54]*tmp[152]+tmp[55]*tmp[151]+tmp[56]*tmp[150]+tmp[57]*tmp[149]+tmp[58]*tmp[148]+tmp[59]*tmp[147]+tmp[60]*tmp[146]+tmp[61]*tmp[145]+tmp[62]*tmp[144]+tmp[63]*tmp[143]+tmp[64]*tmp[142]+tmp[65]*tmp[141]+tmp[66]*tmp[140]+tmp[67]*tmp[139]+tmp[68]*tmp[138]+tmp[69]*tmp[137]+tmp[70]*tmp[136]+tmp[71]*tmp[135]+tmp[72]*tmp[134]+tmp[73]*tmp[133]+tmp[74]*tmp[132]+tmp[75]*tmp[131]+tmp[76]*tmp[130]+tmp[77]*tmp[129]+tmp[78]*tmp[128]+tmp[79]*tmp[127]+tmp[80]*tmp[126]+tmp[81]*tmp[125]+tmp[82]*tmp[124]+tmp[83]*tmp[123]+tmp[84]*tmp[122]+tmp[85]*tmp[121]+tmp[86]*tmp[120]+tmp[87]*tmp[119]+tmp[88]*tmp[118]+tmp[89]*tmp[117]+tmp[90]*tmp[116]+tmp[91]*tmp[115]+tmp[92]*tmp[114]+tmp[93]*tmp[113]+tmp[94]*tmp[112]+tmp[95]*tmp[111]+tmp[96]*tmp[110]+tmp[97]*tmp[109]+tmp[98]*tmp[108]+tmp[99]*tmp[107];
				ans[107]<=tmp[8]*tmp[199]+tmp[9]*tmp[198]+tmp[10]*tmp[197]+tmp[11]*tmp[196]+tmp[12]*tmp[195]+tmp[13]*tmp[194]+tmp[14]*tmp[193]+tmp[15]*tmp[192]+tmp[16]*tmp[191]+tmp[17]*tmp[190]+tmp[18]*tmp[189]+tmp[19]*tmp[188]+tmp[20]*tmp[187]+tmp[21]*tmp[186]+tmp[22]*tmp[185]+tmp[23]*tmp[184]+tmp[24]*tmp[183]+tmp[25]*tmp[182]+tmp[26]*tmp[181]+tmp[27]*tmp[180]+tmp[28]*tmp[179]+tmp[29]*tmp[178]+tmp[30]*tmp[177]+tmp[31]*tmp[176]+tmp[32]*tmp[175]+tmp[33]*tmp[174]+tmp[34]*tmp[173]+tmp[35]*tmp[172]+tmp[36]*tmp[171]+tmp[37]*tmp[170]+tmp[38]*tmp[169]+tmp[39]*tmp[168]+tmp[40]*tmp[167]+tmp[41]*tmp[166]+tmp[42]*tmp[165]+tmp[43]*tmp[164]+tmp[44]*tmp[163]+tmp[45]*tmp[162]+tmp[46]*tmp[161]+tmp[47]*tmp[160]+tmp[48]*tmp[159]+tmp[49]*tmp[158]+tmp[50]*tmp[157]+tmp[51]*tmp[156]+tmp[52]*tmp[155]+tmp[53]*tmp[154]+tmp[54]*tmp[153]+tmp[55]*tmp[152]+tmp[56]*tmp[151]+tmp[57]*tmp[150]+tmp[58]*tmp[149]+tmp[59]*tmp[148]+tmp[60]*tmp[147]+tmp[61]*tmp[146]+tmp[62]*tmp[145]+tmp[63]*tmp[144]+tmp[64]*tmp[143]+tmp[65]*tmp[142]+tmp[66]*tmp[141]+tmp[67]*tmp[140]+tmp[68]*tmp[139]+tmp[69]*tmp[138]+tmp[70]*tmp[137]+tmp[71]*tmp[136]+tmp[72]*tmp[135]+tmp[73]*tmp[134]+tmp[74]*tmp[133]+tmp[75]*tmp[132]+tmp[76]*tmp[131]+tmp[77]*tmp[130]+tmp[78]*tmp[129]+tmp[79]*tmp[128]+tmp[80]*tmp[127]+tmp[81]*tmp[126]+tmp[82]*tmp[125]+tmp[83]*tmp[124]+tmp[84]*tmp[123]+tmp[85]*tmp[122]+tmp[86]*tmp[121]+tmp[87]*tmp[120]+tmp[88]*tmp[119]+tmp[89]*tmp[118]+tmp[90]*tmp[117]+tmp[91]*tmp[116]+tmp[92]*tmp[115]+tmp[93]*tmp[114]+tmp[94]*tmp[113]+tmp[95]*tmp[112]+tmp[96]*tmp[111]+tmp[97]*tmp[110]+tmp[98]*tmp[109]+tmp[99]*tmp[108];
				ans[108]<=tmp[9]*tmp[199]+tmp[10]*tmp[198]+tmp[11]*tmp[197]+tmp[12]*tmp[196]+tmp[13]*tmp[195]+tmp[14]*tmp[194]+tmp[15]*tmp[193]+tmp[16]*tmp[192]+tmp[17]*tmp[191]+tmp[18]*tmp[190]+tmp[19]*tmp[189]+tmp[20]*tmp[188]+tmp[21]*tmp[187]+tmp[22]*tmp[186]+tmp[23]*tmp[185]+tmp[24]*tmp[184]+tmp[25]*tmp[183]+tmp[26]*tmp[182]+tmp[27]*tmp[181]+tmp[28]*tmp[180]+tmp[29]*tmp[179]+tmp[30]*tmp[178]+tmp[31]*tmp[177]+tmp[32]*tmp[176]+tmp[33]*tmp[175]+tmp[34]*tmp[174]+tmp[35]*tmp[173]+tmp[36]*tmp[172]+tmp[37]*tmp[171]+tmp[38]*tmp[170]+tmp[39]*tmp[169]+tmp[40]*tmp[168]+tmp[41]*tmp[167]+tmp[42]*tmp[166]+tmp[43]*tmp[165]+tmp[44]*tmp[164]+tmp[45]*tmp[163]+tmp[46]*tmp[162]+tmp[47]*tmp[161]+tmp[48]*tmp[160]+tmp[49]*tmp[159]+tmp[50]*tmp[158]+tmp[51]*tmp[157]+tmp[52]*tmp[156]+tmp[53]*tmp[155]+tmp[54]*tmp[154]+tmp[55]*tmp[153]+tmp[56]*tmp[152]+tmp[57]*tmp[151]+tmp[58]*tmp[150]+tmp[59]*tmp[149]+tmp[60]*tmp[148]+tmp[61]*tmp[147]+tmp[62]*tmp[146]+tmp[63]*tmp[145]+tmp[64]*tmp[144]+tmp[65]*tmp[143]+tmp[66]*tmp[142]+tmp[67]*tmp[141]+tmp[68]*tmp[140]+tmp[69]*tmp[139]+tmp[70]*tmp[138]+tmp[71]*tmp[137]+tmp[72]*tmp[136]+tmp[73]*tmp[135]+tmp[74]*tmp[134]+tmp[75]*tmp[133]+tmp[76]*tmp[132]+tmp[77]*tmp[131]+tmp[78]*tmp[130]+tmp[79]*tmp[129]+tmp[80]*tmp[128]+tmp[81]*tmp[127]+tmp[82]*tmp[126]+tmp[83]*tmp[125]+tmp[84]*tmp[124]+tmp[85]*tmp[123]+tmp[86]*tmp[122]+tmp[87]*tmp[121]+tmp[88]*tmp[120]+tmp[89]*tmp[119]+tmp[90]*tmp[118]+tmp[91]*tmp[117]+tmp[92]*tmp[116]+tmp[93]*tmp[115]+tmp[94]*tmp[114]+tmp[95]*tmp[113]+tmp[96]*tmp[112]+tmp[97]*tmp[111]+tmp[98]*tmp[110]+tmp[99]*tmp[109];
				ans[109]<=tmp[10]*tmp[199]+tmp[11]*tmp[198]+tmp[12]*tmp[197]+tmp[13]*tmp[196]+tmp[14]*tmp[195]+tmp[15]*tmp[194]+tmp[16]*tmp[193]+tmp[17]*tmp[192]+tmp[18]*tmp[191]+tmp[19]*tmp[190]+tmp[20]*tmp[189]+tmp[21]*tmp[188]+tmp[22]*tmp[187]+tmp[23]*tmp[186]+tmp[24]*tmp[185]+tmp[25]*tmp[184]+tmp[26]*tmp[183]+tmp[27]*tmp[182]+tmp[28]*tmp[181]+tmp[29]*tmp[180]+tmp[30]*tmp[179]+tmp[31]*tmp[178]+tmp[32]*tmp[177]+tmp[33]*tmp[176]+tmp[34]*tmp[175]+tmp[35]*tmp[174]+tmp[36]*tmp[173]+tmp[37]*tmp[172]+tmp[38]*tmp[171]+tmp[39]*tmp[170]+tmp[40]*tmp[169]+tmp[41]*tmp[168]+tmp[42]*tmp[167]+tmp[43]*tmp[166]+tmp[44]*tmp[165]+tmp[45]*tmp[164]+tmp[46]*tmp[163]+tmp[47]*tmp[162]+tmp[48]*tmp[161]+tmp[49]*tmp[160]+tmp[50]*tmp[159]+tmp[51]*tmp[158]+tmp[52]*tmp[157]+tmp[53]*tmp[156]+tmp[54]*tmp[155]+tmp[55]*tmp[154]+tmp[56]*tmp[153]+tmp[57]*tmp[152]+tmp[58]*tmp[151]+tmp[59]*tmp[150]+tmp[60]*tmp[149]+tmp[61]*tmp[148]+tmp[62]*tmp[147]+tmp[63]*tmp[146]+tmp[64]*tmp[145]+tmp[65]*tmp[144]+tmp[66]*tmp[143]+tmp[67]*tmp[142]+tmp[68]*tmp[141]+tmp[69]*tmp[140]+tmp[70]*tmp[139]+tmp[71]*tmp[138]+tmp[72]*tmp[137]+tmp[73]*tmp[136]+tmp[74]*tmp[135]+tmp[75]*tmp[134]+tmp[76]*tmp[133]+tmp[77]*tmp[132]+tmp[78]*tmp[131]+tmp[79]*tmp[130]+tmp[80]*tmp[129]+tmp[81]*tmp[128]+tmp[82]*tmp[127]+tmp[83]*tmp[126]+tmp[84]*tmp[125]+tmp[85]*tmp[124]+tmp[86]*tmp[123]+tmp[87]*tmp[122]+tmp[88]*tmp[121]+tmp[89]*tmp[120]+tmp[90]*tmp[119]+tmp[91]*tmp[118]+tmp[92]*tmp[117]+tmp[93]*tmp[116]+tmp[94]*tmp[115]+tmp[95]*tmp[114]+tmp[96]*tmp[113]+tmp[97]*tmp[112]+tmp[98]*tmp[111]+tmp[99]*tmp[110];
				ans[110]<=tmp[11]*tmp[199]+tmp[12]*tmp[198]+tmp[13]*tmp[197]+tmp[14]*tmp[196]+tmp[15]*tmp[195]+tmp[16]*tmp[194]+tmp[17]*tmp[193]+tmp[18]*tmp[192]+tmp[19]*tmp[191]+tmp[20]*tmp[190]+tmp[21]*tmp[189]+tmp[22]*tmp[188]+tmp[23]*tmp[187]+tmp[24]*tmp[186]+tmp[25]*tmp[185]+tmp[26]*tmp[184]+tmp[27]*tmp[183]+tmp[28]*tmp[182]+tmp[29]*tmp[181]+tmp[30]*tmp[180]+tmp[31]*tmp[179]+tmp[32]*tmp[178]+tmp[33]*tmp[177]+tmp[34]*tmp[176]+tmp[35]*tmp[175]+tmp[36]*tmp[174]+tmp[37]*tmp[173]+tmp[38]*tmp[172]+tmp[39]*tmp[171]+tmp[40]*tmp[170]+tmp[41]*tmp[169]+tmp[42]*tmp[168]+tmp[43]*tmp[167]+tmp[44]*tmp[166]+tmp[45]*tmp[165]+tmp[46]*tmp[164]+tmp[47]*tmp[163]+tmp[48]*tmp[162]+tmp[49]*tmp[161]+tmp[50]*tmp[160]+tmp[51]*tmp[159]+tmp[52]*tmp[158]+tmp[53]*tmp[157]+tmp[54]*tmp[156]+tmp[55]*tmp[155]+tmp[56]*tmp[154]+tmp[57]*tmp[153]+tmp[58]*tmp[152]+tmp[59]*tmp[151]+tmp[60]*tmp[150]+tmp[61]*tmp[149]+tmp[62]*tmp[148]+tmp[63]*tmp[147]+tmp[64]*tmp[146]+tmp[65]*tmp[145]+tmp[66]*tmp[144]+tmp[67]*tmp[143]+tmp[68]*tmp[142]+tmp[69]*tmp[141]+tmp[70]*tmp[140]+tmp[71]*tmp[139]+tmp[72]*tmp[138]+tmp[73]*tmp[137]+tmp[74]*tmp[136]+tmp[75]*tmp[135]+tmp[76]*tmp[134]+tmp[77]*tmp[133]+tmp[78]*tmp[132]+tmp[79]*tmp[131]+tmp[80]*tmp[130]+tmp[81]*tmp[129]+tmp[82]*tmp[128]+tmp[83]*tmp[127]+tmp[84]*tmp[126]+tmp[85]*tmp[125]+tmp[86]*tmp[124]+tmp[87]*tmp[123]+tmp[88]*tmp[122]+tmp[89]*tmp[121]+tmp[90]*tmp[120]+tmp[91]*tmp[119]+tmp[92]*tmp[118]+tmp[93]*tmp[117]+tmp[94]*tmp[116]+tmp[95]*tmp[115]+tmp[96]*tmp[114]+tmp[97]*tmp[113]+tmp[98]*tmp[112]+tmp[99]*tmp[111];
				ans[111]<=tmp[12]*tmp[199]+tmp[13]*tmp[198]+tmp[14]*tmp[197]+tmp[15]*tmp[196]+tmp[16]*tmp[195]+tmp[17]*tmp[194]+tmp[18]*tmp[193]+tmp[19]*tmp[192]+tmp[20]*tmp[191]+tmp[21]*tmp[190]+tmp[22]*tmp[189]+tmp[23]*tmp[188]+tmp[24]*tmp[187]+tmp[25]*tmp[186]+tmp[26]*tmp[185]+tmp[27]*tmp[184]+tmp[28]*tmp[183]+tmp[29]*tmp[182]+tmp[30]*tmp[181]+tmp[31]*tmp[180]+tmp[32]*tmp[179]+tmp[33]*tmp[178]+tmp[34]*tmp[177]+tmp[35]*tmp[176]+tmp[36]*tmp[175]+tmp[37]*tmp[174]+tmp[38]*tmp[173]+tmp[39]*tmp[172]+tmp[40]*tmp[171]+tmp[41]*tmp[170]+tmp[42]*tmp[169]+tmp[43]*tmp[168]+tmp[44]*tmp[167]+tmp[45]*tmp[166]+tmp[46]*tmp[165]+tmp[47]*tmp[164]+tmp[48]*tmp[163]+tmp[49]*tmp[162]+tmp[50]*tmp[161]+tmp[51]*tmp[160]+tmp[52]*tmp[159]+tmp[53]*tmp[158]+tmp[54]*tmp[157]+tmp[55]*tmp[156]+tmp[56]*tmp[155]+tmp[57]*tmp[154]+tmp[58]*tmp[153]+tmp[59]*tmp[152]+tmp[60]*tmp[151]+tmp[61]*tmp[150]+tmp[62]*tmp[149]+tmp[63]*tmp[148]+tmp[64]*tmp[147]+tmp[65]*tmp[146]+tmp[66]*tmp[145]+tmp[67]*tmp[144]+tmp[68]*tmp[143]+tmp[69]*tmp[142]+tmp[70]*tmp[141]+tmp[71]*tmp[140]+tmp[72]*tmp[139]+tmp[73]*tmp[138]+tmp[74]*tmp[137]+tmp[75]*tmp[136]+tmp[76]*tmp[135]+tmp[77]*tmp[134]+tmp[78]*tmp[133]+tmp[79]*tmp[132]+tmp[80]*tmp[131]+tmp[81]*tmp[130]+tmp[82]*tmp[129]+tmp[83]*tmp[128]+tmp[84]*tmp[127]+tmp[85]*tmp[126]+tmp[86]*tmp[125]+tmp[87]*tmp[124]+tmp[88]*tmp[123]+tmp[89]*tmp[122]+tmp[90]*tmp[121]+tmp[91]*tmp[120]+tmp[92]*tmp[119]+tmp[93]*tmp[118]+tmp[94]*tmp[117]+tmp[95]*tmp[116]+tmp[96]*tmp[115]+tmp[97]*tmp[114]+tmp[98]*tmp[113]+tmp[99]*tmp[112];
				ans[112]<=tmp[13]*tmp[199]+tmp[14]*tmp[198]+tmp[15]*tmp[197]+tmp[16]*tmp[196]+tmp[17]*tmp[195]+tmp[18]*tmp[194]+tmp[19]*tmp[193]+tmp[20]*tmp[192]+tmp[21]*tmp[191]+tmp[22]*tmp[190]+tmp[23]*tmp[189]+tmp[24]*tmp[188]+tmp[25]*tmp[187]+tmp[26]*tmp[186]+tmp[27]*tmp[185]+tmp[28]*tmp[184]+tmp[29]*tmp[183]+tmp[30]*tmp[182]+tmp[31]*tmp[181]+tmp[32]*tmp[180]+tmp[33]*tmp[179]+tmp[34]*tmp[178]+tmp[35]*tmp[177]+tmp[36]*tmp[176]+tmp[37]*tmp[175]+tmp[38]*tmp[174]+tmp[39]*tmp[173]+tmp[40]*tmp[172]+tmp[41]*tmp[171]+tmp[42]*tmp[170]+tmp[43]*tmp[169]+tmp[44]*tmp[168]+tmp[45]*tmp[167]+tmp[46]*tmp[166]+tmp[47]*tmp[165]+tmp[48]*tmp[164]+tmp[49]*tmp[163]+tmp[50]*tmp[162]+tmp[51]*tmp[161]+tmp[52]*tmp[160]+tmp[53]*tmp[159]+tmp[54]*tmp[158]+tmp[55]*tmp[157]+tmp[56]*tmp[156]+tmp[57]*tmp[155]+tmp[58]*tmp[154]+tmp[59]*tmp[153]+tmp[60]*tmp[152]+tmp[61]*tmp[151]+tmp[62]*tmp[150]+tmp[63]*tmp[149]+tmp[64]*tmp[148]+tmp[65]*tmp[147]+tmp[66]*tmp[146]+tmp[67]*tmp[145]+tmp[68]*tmp[144]+tmp[69]*tmp[143]+tmp[70]*tmp[142]+tmp[71]*tmp[141]+tmp[72]*tmp[140]+tmp[73]*tmp[139]+tmp[74]*tmp[138]+tmp[75]*tmp[137]+tmp[76]*tmp[136]+tmp[77]*tmp[135]+tmp[78]*tmp[134]+tmp[79]*tmp[133]+tmp[80]*tmp[132]+tmp[81]*tmp[131]+tmp[82]*tmp[130]+tmp[83]*tmp[129]+tmp[84]*tmp[128]+tmp[85]*tmp[127]+tmp[86]*tmp[126]+tmp[87]*tmp[125]+tmp[88]*tmp[124]+tmp[89]*tmp[123]+tmp[90]*tmp[122]+tmp[91]*tmp[121]+tmp[92]*tmp[120]+tmp[93]*tmp[119]+tmp[94]*tmp[118]+tmp[95]*tmp[117]+tmp[96]*tmp[116]+tmp[97]*tmp[115]+tmp[98]*tmp[114]+tmp[99]*tmp[113];
				ans[113]<=tmp[14]*tmp[199]+tmp[15]*tmp[198]+tmp[16]*tmp[197]+tmp[17]*tmp[196]+tmp[18]*tmp[195]+tmp[19]*tmp[194]+tmp[20]*tmp[193]+tmp[21]*tmp[192]+tmp[22]*tmp[191]+tmp[23]*tmp[190]+tmp[24]*tmp[189]+tmp[25]*tmp[188]+tmp[26]*tmp[187]+tmp[27]*tmp[186]+tmp[28]*tmp[185]+tmp[29]*tmp[184]+tmp[30]*tmp[183]+tmp[31]*tmp[182]+tmp[32]*tmp[181]+tmp[33]*tmp[180]+tmp[34]*tmp[179]+tmp[35]*tmp[178]+tmp[36]*tmp[177]+tmp[37]*tmp[176]+tmp[38]*tmp[175]+tmp[39]*tmp[174]+tmp[40]*tmp[173]+tmp[41]*tmp[172]+tmp[42]*tmp[171]+tmp[43]*tmp[170]+tmp[44]*tmp[169]+tmp[45]*tmp[168]+tmp[46]*tmp[167]+tmp[47]*tmp[166]+tmp[48]*tmp[165]+tmp[49]*tmp[164]+tmp[50]*tmp[163]+tmp[51]*tmp[162]+tmp[52]*tmp[161]+tmp[53]*tmp[160]+tmp[54]*tmp[159]+tmp[55]*tmp[158]+tmp[56]*tmp[157]+tmp[57]*tmp[156]+tmp[58]*tmp[155]+tmp[59]*tmp[154]+tmp[60]*tmp[153]+tmp[61]*tmp[152]+tmp[62]*tmp[151]+tmp[63]*tmp[150]+tmp[64]*tmp[149]+tmp[65]*tmp[148]+tmp[66]*tmp[147]+tmp[67]*tmp[146]+tmp[68]*tmp[145]+tmp[69]*tmp[144]+tmp[70]*tmp[143]+tmp[71]*tmp[142]+tmp[72]*tmp[141]+tmp[73]*tmp[140]+tmp[74]*tmp[139]+tmp[75]*tmp[138]+tmp[76]*tmp[137]+tmp[77]*tmp[136]+tmp[78]*tmp[135]+tmp[79]*tmp[134]+tmp[80]*tmp[133]+tmp[81]*tmp[132]+tmp[82]*tmp[131]+tmp[83]*tmp[130]+tmp[84]*tmp[129]+tmp[85]*tmp[128]+tmp[86]*tmp[127]+tmp[87]*tmp[126]+tmp[88]*tmp[125]+tmp[89]*tmp[124]+tmp[90]*tmp[123]+tmp[91]*tmp[122]+tmp[92]*tmp[121]+tmp[93]*tmp[120]+tmp[94]*tmp[119]+tmp[95]*tmp[118]+tmp[96]*tmp[117]+tmp[97]*tmp[116]+tmp[98]*tmp[115]+tmp[99]*tmp[114];
				ans[114]<=tmp[15]*tmp[199]+tmp[16]*tmp[198]+tmp[17]*tmp[197]+tmp[18]*tmp[196]+tmp[19]*tmp[195]+tmp[20]*tmp[194]+tmp[21]*tmp[193]+tmp[22]*tmp[192]+tmp[23]*tmp[191]+tmp[24]*tmp[190]+tmp[25]*tmp[189]+tmp[26]*tmp[188]+tmp[27]*tmp[187]+tmp[28]*tmp[186]+tmp[29]*tmp[185]+tmp[30]*tmp[184]+tmp[31]*tmp[183]+tmp[32]*tmp[182]+tmp[33]*tmp[181]+tmp[34]*tmp[180]+tmp[35]*tmp[179]+tmp[36]*tmp[178]+tmp[37]*tmp[177]+tmp[38]*tmp[176]+tmp[39]*tmp[175]+tmp[40]*tmp[174]+tmp[41]*tmp[173]+tmp[42]*tmp[172]+tmp[43]*tmp[171]+tmp[44]*tmp[170]+tmp[45]*tmp[169]+tmp[46]*tmp[168]+tmp[47]*tmp[167]+tmp[48]*tmp[166]+tmp[49]*tmp[165]+tmp[50]*tmp[164]+tmp[51]*tmp[163]+tmp[52]*tmp[162]+tmp[53]*tmp[161]+tmp[54]*tmp[160]+tmp[55]*tmp[159]+tmp[56]*tmp[158]+tmp[57]*tmp[157]+tmp[58]*tmp[156]+tmp[59]*tmp[155]+tmp[60]*tmp[154]+tmp[61]*tmp[153]+tmp[62]*tmp[152]+tmp[63]*tmp[151]+tmp[64]*tmp[150]+tmp[65]*tmp[149]+tmp[66]*tmp[148]+tmp[67]*tmp[147]+tmp[68]*tmp[146]+tmp[69]*tmp[145]+tmp[70]*tmp[144]+tmp[71]*tmp[143]+tmp[72]*tmp[142]+tmp[73]*tmp[141]+tmp[74]*tmp[140]+tmp[75]*tmp[139]+tmp[76]*tmp[138]+tmp[77]*tmp[137]+tmp[78]*tmp[136]+tmp[79]*tmp[135]+tmp[80]*tmp[134]+tmp[81]*tmp[133]+tmp[82]*tmp[132]+tmp[83]*tmp[131]+tmp[84]*tmp[130]+tmp[85]*tmp[129]+tmp[86]*tmp[128]+tmp[87]*tmp[127]+tmp[88]*tmp[126]+tmp[89]*tmp[125]+tmp[90]*tmp[124]+tmp[91]*tmp[123]+tmp[92]*tmp[122]+tmp[93]*tmp[121]+tmp[94]*tmp[120]+tmp[95]*tmp[119]+tmp[96]*tmp[118]+tmp[97]*tmp[117]+tmp[98]*tmp[116]+tmp[99]*tmp[115];
				ans[115]<=tmp[16]*tmp[199]+tmp[17]*tmp[198]+tmp[18]*tmp[197]+tmp[19]*tmp[196]+tmp[20]*tmp[195]+tmp[21]*tmp[194]+tmp[22]*tmp[193]+tmp[23]*tmp[192]+tmp[24]*tmp[191]+tmp[25]*tmp[190]+tmp[26]*tmp[189]+tmp[27]*tmp[188]+tmp[28]*tmp[187]+tmp[29]*tmp[186]+tmp[30]*tmp[185]+tmp[31]*tmp[184]+tmp[32]*tmp[183]+tmp[33]*tmp[182]+tmp[34]*tmp[181]+tmp[35]*tmp[180]+tmp[36]*tmp[179]+tmp[37]*tmp[178]+tmp[38]*tmp[177]+tmp[39]*tmp[176]+tmp[40]*tmp[175]+tmp[41]*tmp[174]+tmp[42]*tmp[173]+tmp[43]*tmp[172]+tmp[44]*tmp[171]+tmp[45]*tmp[170]+tmp[46]*tmp[169]+tmp[47]*tmp[168]+tmp[48]*tmp[167]+tmp[49]*tmp[166]+tmp[50]*tmp[165]+tmp[51]*tmp[164]+tmp[52]*tmp[163]+tmp[53]*tmp[162]+tmp[54]*tmp[161]+tmp[55]*tmp[160]+tmp[56]*tmp[159]+tmp[57]*tmp[158]+tmp[58]*tmp[157]+tmp[59]*tmp[156]+tmp[60]*tmp[155]+tmp[61]*tmp[154]+tmp[62]*tmp[153]+tmp[63]*tmp[152]+tmp[64]*tmp[151]+tmp[65]*tmp[150]+tmp[66]*tmp[149]+tmp[67]*tmp[148]+tmp[68]*tmp[147]+tmp[69]*tmp[146]+tmp[70]*tmp[145]+tmp[71]*tmp[144]+tmp[72]*tmp[143]+tmp[73]*tmp[142]+tmp[74]*tmp[141]+tmp[75]*tmp[140]+tmp[76]*tmp[139]+tmp[77]*tmp[138]+tmp[78]*tmp[137]+tmp[79]*tmp[136]+tmp[80]*tmp[135]+tmp[81]*tmp[134]+tmp[82]*tmp[133]+tmp[83]*tmp[132]+tmp[84]*tmp[131]+tmp[85]*tmp[130]+tmp[86]*tmp[129]+tmp[87]*tmp[128]+tmp[88]*tmp[127]+tmp[89]*tmp[126]+tmp[90]*tmp[125]+tmp[91]*tmp[124]+tmp[92]*tmp[123]+tmp[93]*tmp[122]+tmp[94]*tmp[121]+tmp[95]*tmp[120]+tmp[96]*tmp[119]+tmp[97]*tmp[118]+tmp[98]*tmp[117]+tmp[99]*tmp[116];
				ans[116]<=tmp[17]*tmp[199]+tmp[18]*tmp[198]+tmp[19]*tmp[197]+tmp[20]*tmp[196]+tmp[21]*tmp[195]+tmp[22]*tmp[194]+tmp[23]*tmp[193]+tmp[24]*tmp[192]+tmp[25]*tmp[191]+tmp[26]*tmp[190]+tmp[27]*tmp[189]+tmp[28]*tmp[188]+tmp[29]*tmp[187]+tmp[30]*tmp[186]+tmp[31]*tmp[185]+tmp[32]*tmp[184]+tmp[33]*tmp[183]+tmp[34]*tmp[182]+tmp[35]*tmp[181]+tmp[36]*tmp[180]+tmp[37]*tmp[179]+tmp[38]*tmp[178]+tmp[39]*tmp[177]+tmp[40]*tmp[176]+tmp[41]*tmp[175]+tmp[42]*tmp[174]+tmp[43]*tmp[173]+tmp[44]*tmp[172]+tmp[45]*tmp[171]+tmp[46]*tmp[170]+tmp[47]*tmp[169]+tmp[48]*tmp[168]+tmp[49]*tmp[167]+tmp[50]*tmp[166]+tmp[51]*tmp[165]+tmp[52]*tmp[164]+tmp[53]*tmp[163]+tmp[54]*tmp[162]+tmp[55]*tmp[161]+tmp[56]*tmp[160]+tmp[57]*tmp[159]+tmp[58]*tmp[158]+tmp[59]*tmp[157]+tmp[60]*tmp[156]+tmp[61]*tmp[155]+tmp[62]*tmp[154]+tmp[63]*tmp[153]+tmp[64]*tmp[152]+tmp[65]*tmp[151]+tmp[66]*tmp[150]+tmp[67]*tmp[149]+tmp[68]*tmp[148]+tmp[69]*tmp[147]+tmp[70]*tmp[146]+tmp[71]*tmp[145]+tmp[72]*tmp[144]+tmp[73]*tmp[143]+tmp[74]*tmp[142]+tmp[75]*tmp[141]+tmp[76]*tmp[140]+tmp[77]*tmp[139]+tmp[78]*tmp[138]+tmp[79]*tmp[137]+tmp[80]*tmp[136]+tmp[81]*tmp[135]+tmp[82]*tmp[134]+tmp[83]*tmp[133]+tmp[84]*tmp[132]+tmp[85]*tmp[131]+tmp[86]*tmp[130]+tmp[87]*tmp[129]+tmp[88]*tmp[128]+tmp[89]*tmp[127]+tmp[90]*tmp[126]+tmp[91]*tmp[125]+tmp[92]*tmp[124]+tmp[93]*tmp[123]+tmp[94]*tmp[122]+tmp[95]*tmp[121]+tmp[96]*tmp[120]+tmp[97]*tmp[119]+tmp[98]*tmp[118]+tmp[99]*tmp[117];
				ans[117]<=tmp[18]*tmp[199]+tmp[19]*tmp[198]+tmp[20]*tmp[197]+tmp[21]*tmp[196]+tmp[22]*tmp[195]+tmp[23]*tmp[194]+tmp[24]*tmp[193]+tmp[25]*tmp[192]+tmp[26]*tmp[191]+tmp[27]*tmp[190]+tmp[28]*tmp[189]+tmp[29]*tmp[188]+tmp[30]*tmp[187]+tmp[31]*tmp[186]+tmp[32]*tmp[185]+tmp[33]*tmp[184]+tmp[34]*tmp[183]+tmp[35]*tmp[182]+tmp[36]*tmp[181]+tmp[37]*tmp[180]+tmp[38]*tmp[179]+tmp[39]*tmp[178]+tmp[40]*tmp[177]+tmp[41]*tmp[176]+tmp[42]*tmp[175]+tmp[43]*tmp[174]+tmp[44]*tmp[173]+tmp[45]*tmp[172]+tmp[46]*tmp[171]+tmp[47]*tmp[170]+tmp[48]*tmp[169]+tmp[49]*tmp[168]+tmp[50]*tmp[167]+tmp[51]*tmp[166]+tmp[52]*tmp[165]+tmp[53]*tmp[164]+tmp[54]*tmp[163]+tmp[55]*tmp[162]+tmp[56]*tmp[161]+tmp[57]*tmp[160]+tmp[58]*tmp[159]+tmp[59]*tmp[158]+tmp[60]*tmp[157]+tmp[61]*tmp[156]+tmp[62]*tmp[155]+tmp[63]*tmp[154]+tmp[64]*tmp[153]+tmp[65]*tmp[152]+tmp[66]*tmp[151]+tmp[67]*tmp[150]+tmp[68]*tmp[149]+tmp[69]*tmp[148]+tmp[70]*tmp[147]+tmp[71]*tmp[146]+tmp[72]*tmp[145]+tmp[73]*tmp[144]+tmp[74]*tmp[143]+tmp[75]*tmp[142]+tmp[76]*tmp[141]+tmp[77]*tmp[140]+tmp[78]*tmp[139]+tmp[79]*tmp[138]+tmp[80]*tmp[137]+tmp[81]*tmp[136]+tmp[82]*tmp[135]+tmp[83]*tmp[134]+tmp[84]*tmp[133]+tmp[85]*tmp[132]+tmp[86]*tmp[131]+tmp[87]*tmp[130]+tmp[88]*tmp[129]+tmp[89]*tmp[128]+tmp[90]*tmp[127]+tmp[91]*tmp[126]+tmp[92]*tmp[125]+tmp[93]*tmp[124]+tmp[94]*tmp[123]+tmp[95]*tmp[122]+tmp[96]*tmp[121]+tmp[97]*tmp[120]+tmp[98]*tmp[119]+tmp[99]*tmp[118];
				ans[118]<=tmp[19]*tmp[199]+tmp[20]*tmp[198]+tmp[21]*tmp[197]+tmp[22]*tmp[196]+tmp[23]*tmp[195]+tmp[24]*tmp[194]+tmp[25]*tmp[193]+tmp[26]*tmp[192]+tmp[27]*tmp[191]+tmp[28]*tmp[190]+tmp[29]*tmp[189]+tmp[30]*tmp[188]+tmp[31]*tmp[187]+tmp[32]*tmp[186]+tmp[33]*tmp[185]+tmp[34]*tmp[184]+tmp[35]*tmp[183]+tmp[36]*tmp[182]+tmp[37]*tmp[181]+tmp[38]*tmp[180]+tmp[39]*tmp[179]+tmp[40]*tmp[178]+tmp[41]*tmp[177]+tmp[42]*tmp[176]+tmp[43]*tmp[175]+tmp[44]*tmp[174]+tmp[45]*tmp[173]+tmp[46]*tmp[172]+tmp[47]*tmp[171]+tmp[48]*tmp[170]+tmp[49]*tmp[169]+tmp[50]*tmp[168]+tmp[51]*tmp[167]+tmp[52]*tmp[166]+tmp[53]*tmp[165]+tmp[54]*tmp[164]+tmp[55]*tmp[163]+tmp[56]*tmp[162]+tmp[57]*tmp[161]+tmp[58]*tmp[160]+tmp[59]*tmp[159]+tmp[60]*tmp[158]+tmp[61]*tmp[157]+tmp[62]*tmp[156]+tmp[63]*tmp[155]+tmp[64]*tmp[154]+tmp[65]*tmp[153]+tmp[66]*tmp[152]+tmp[67]*tmp[151]+tmp[68]*tmp[150]+tmp[69]*tmp[149]+tmp[70]*tmp[148]+tmp[71]*tmp[147]+tmp[72]*tmp[146]+tmp[73]*tmp[145]+tmp[74]*tmp[144]+tmp[75]*tmp[143]+tmp[76]*tmp[142]+tmp[77]*tmp[141]+tmp[78]*tmp[140]+tmp[79]*tmp[139]+tmp[80]*tmp[138]+tmp[81]*tmp[137]+tmp[82]*tmp[136]+tmp[83]*tmp[135]+tmp[84]*tmp[134]+tmp[85]*tmp[133]+tmp[86]*tmp[132]+tmp[87]*tmp[131]+tmp[88]*tmp[130]+tmp[89]*tmp[129]+tmp[90]*tmp[128]+tmp[91]*tmp[127]+tmp[92]*tmp[126]+tmp[93]*tmp[125]+tmp[94]*tmp[124]+tmp[95]*tmp[123]+tmp[96]*tmp[122]+tmp[97]*tmp[121]+tmp[98]*tmp[120]+tmp[99]*tmp[119];
				ans[119]<=tmp[20]*tmp[199]+tmp[21]*tmp[198]+tmp[22]*tmp[197]+tmp[23]*tmp[196]+tmp[24]*tmp[195]+tmp[25]*tmp[194]+tmp[26]*tmp[193]+tmp[27]*tmp[192]+tmp[28]*tmp[191]+tmp[29]*tmp[190]+tmp[30]*tmp[189]+tmp[31]*tmp[188]+tmp[32]*tmp[187]+tmp[33]*tmp[186]+tmp[34]*tmp[185]+tmp[35]*tmp[184]+tmp[36]*tmp[183]+tmp[37]*tmp[182]+tmp[38]*tmp[181]+tmp[39]*tmp[180]+tmp[40]*tmp[179]+tmp[41]*tmp[178]+tmp[42]*tmp[177]+tmp[43]*tmp[176]+tmp[44]*tmp[175]+tmp[45]*tmp[174]+tmp[46]*tmp[173]+tmp[47]*tmp[172]+tmp[48]*tmp[171]+tmp[49]*tmp[170]+tmp[50]*tmp[169]+tmp[51]*tmp[168]+tmp[52]*tmp[167]+tmp[53]*tmp[166]+tmp[54]*tmp[165]+tmp[55]*tmp[164]+tmp[56]*tmp[163]+tmp[57]*tmp[162]+tmp[58]*tmp[161]+tmp[59]*tmp[160]+tmp[60]*tmp[159]+tmp[61]*tmp[158]+tmp[62]*tmp[157]+tmp[63]*tmp[156]+tmp[64]*tmp[155]+tmp[65]*tmp[154]+tmp[66]*tmp[153]+tmp[67]*tmp[152]+tmp[68]*tmp[151]+tmp[69]*tmp[150]+tmp[70]*tmp[149]+tmp[71]*tmp[148]+tmp[72]*tmp[147]+tmp[73]*tmp[146]+tmp[74]*tmp[145]+tmp[75]*tmp[144]+tmp[76]*tmp[143]+tmp[77]*tmp[142]+tmp[78]*tmp[141]+tmp[79]*tmp[140]+tmp[80]*tmp[139]+tmp[81]*tmp[138]+tmp[82]*tmp[137]+tmp[83]*tmp[136]+tmp[84]*tmp[135]+tmp[85]*tmp[134]+tmp[86]*tmp[133]+tmp[87]*tmp[132]+tmp[88]*tmp[131]+tmp[89]*tmp[130]+tmp[90]*tmp[129]+tmp[91]*tmp[128]+tmp[92]*tmp[127]+tmp[93]*tmp[126]+tmp[94]*tmp[125]+tmp[95]*tmp[124]+tmp[96]*tmp[123]+tmp[97]*tmp[122]+tmp[98]*tmp[121]+tmp[99]*tmp[120];
				ans[120]<=tmp[21]*tmp[199]+tmp[22]*tmp[198]+tmp[23]*tmp[197]+tmp[24]*tmp[196]+tmp[25]*tmp[195]+tmp[26]*tmp[194]+tmp[27]*tmp[193]+tmp[28]*tmp[192]+tmp[29]*tmp[191]+tmp[30]*tmp[190]+tmp[31]*tmp[189]+tmp[32]*tmp[188]+tmp[33]*tmp[187]+tmp[34]*tmp[186]+tmp[35]*tmp[185]+tmp[36]*tmp[184]+tmp[37]*tmp[183]+tmp[38]*tmp[182]+tmp[39]*tmp[181]+tmp[40]*tmp[180]+tmp[41]*tmp[179]+tmp[42]*tmp[178]+tmp[43]*tmp[177]+tmp[44]*tmp[176]+tmp[45]*tmp[175]+tmp[46]*tmp[174]+tmp[47]*tmp[173]+tmp[48]*tmp[172]+tmp[49]*tmp[171]+tmp[50]*tmp[170]+tmp[51]*tmp[169]+tmp[52]*tmp[168]+tmp[53]*tmp[167]+tmp[54]*tmp[166]+tmp[55]*tmp[165]+tmp[56]*tmp[164]+tmp[57]*tmp[163]+tmp[58]*tmp[162]+tmp[59]*tmp[161]+tmp[60]*tmp[160]+tmp[61]*tmp[159]+tmp[62]*tmp[158]+tmp[63]*tmp[157]+tmp[64]*tmp[156]+tmp[65]*tmp[155]+tmp[66]*tmp[154]+tmp[67]*tmp[153]+tmp[68]*tmp[152]+tmp[69]*tmp[151]+tmp[70]*tmp[150]+tmp[71]*tmp[149]+tmp[72]*tmp[148]+tmp[73]*tmp[147]+tmp[74]*tmp[146]+tmp[75]*tmp[145]+tmp[76]*tmp[144]+tmp[77]*tmp[143]+tmp[78]*tmp[142]+tmp[79]*tmp[141]+tmp[80]*tmp[140]+tmp[81]*tmp[139]+tmp[82]*tmp[138]+tmp[83]*tmp[137]+tmp[84]*tmp[136]+tmp[85]*tmp[135]+tmp[86]*tmp[134]+tmp[87]*tmp[133]+tmp[88]*tmp[132]+tmp[89]*tmp[131]+tmp[90]*tmp[130]+tmp[91]*tmp[129]+tmp[92]*tmp[128]+tmp[93]*tmp[127]+tmp[94]*tmp[126]+tmp[95]*tmp[125]+tmp[96]*tmp[124]+tmp[97]*tmp[123]+tmp[98]*tmp[122]+tmp[99]*tmp[121];
				ans[121]<=tmp[22]*tmp[199]+tmp[23]*tmp[198]+tmp[24]*tmp[197]+tmp[25]*tmp[196]+tmp[26]*tmp[195]+tmp[27]*tmp[194]+tmp[28]*tmp[193]+tmp[29]*tmp[192]+tmp[30]*tmp[191]+tmp[31]*tmp[190]+tmp[32]*tmp[189]+tmp[33]*tmp[188]+tmp[34]*tmp[187]+tmp[35]*tmp[186]+tmp[36]*tmp[185]+tmp[37]*tmp[184]+tmp[38]*tmp[183]+tmp[39]*tmp[182]+tmp[40]*tmp[181]+tmp[41]*tmp[180]+tmp[42]*tmp[179]+tmp[43]*tmp[178]+tmp[44]*tmp[177]+tmp[45]*tmp[176]+tmp[46]*tmp[175]+tmp[47]*tmp[174]+tmp[48]*tmp[173]+tmp[49]*tmp[172]+tmp[50]*tmp[171]+tmp[51]*tmp[170]+tmp[52]*tmp[169]+tmp[53]*tmp[168]+tmp[54]*tmp[167]+tmp[55]*tmp[166]+tmp[56]*tmp[165]+tmp[57]*tmp[164]+tmp[58]*tmp[163]+tmp[59]*tmp[162]+tmp[60]*tmp[161]+tmp[61]*tmp[160]+tmp[62]*tmp[159]+tmp[63]*tmp[158]+tmp[64]*tmp[157]+tmp[65]*tmp[156]+tmp[66]*tmp[155]+tmp[67]*tmp[154]+tmp[68]*tmp[153]+tmp[69]*tmp[152]+tmp[70]*tmp[151]+tmp[71]*tmp[150]+tmp[72]*tmp[149]+tmp[73]*tmp[148]+tmp[74]*tmp[147]+tmp[75]*tmp[146]+tmp[76]*tmp[145]+tmp[77]*tmp[144]+tmp[78]*tmp[143]+tmp[79]*tmp[142]+tmp[80]*tmp[141]+tmp[81]*tmp[140]+tmp[82]*tmp[139]+tmp[83]*tmp[138]+tmp[84]*tmp[137]+tmp[85]*tmp[136]+tmp[86]*tmp[135]+tmp[87]*tmp[134]+tmp[88]*tmp[133]+tmp[89]*tmp[132]+tmp[90]*tmp[131]+tmp[91]*tmp[130]+tmp[92]*tmp[129]+tmp[93]*tmp[128]+tmp[94]*tmp[127]+tmp[95]*tmp[126]+tmp[96]*tmp[125]+tmp[97]*tmp[124]+tmp[98]*tmp[123]+tmp[99]*tmp[122];
				ans[122]<=tmp[23]*tmp[199]+tmp[24]*tmp[198]+tmp[25]*tmp[197]+tmp[26]*tmp[196]+tmp[27]*tmp[195]+tmp[28]*tmp[194]+tmp[29]*tmp[193]+tmp[30]*tmp[192]+tmp[31]*tmp[191]+tmp[32]*tmp[190]+tmp[33]*tmp[189]+tmp[34]*tmp[188]+tmp[35]*tmp[187]+tmp[36]*tmp[186]+tmp[37]*tmp[185]+tmp[38]*tmp[184]+tmp[39]*tmp[183]+tmp[40]*tmp[182]+tmp[41]*tmp[181]+tmp[42]*tmp[180]+tmp[43]*tmp[179]+tmp[44]*tmp[178]+tmp[45]*tmp[177]+tmp[46]*tmp[176]+tmp[47]*tmp[175]+tmp[48]*tmp[174]+tmp[49]*tmp[173]+tmp[50]*tmp[172]+tmp[51]*tmp[171]+tmp[52]*tmp[170]+tmp[53]*tmp[169]+tmp[54]*tmp[168]+tmp[55]*tmp[167]+tmp[56]*tmp[166]+tmp[57]*tmp[165]+tmp[58]*tmp[164]+tmp[59]*tmp[163]+tmp[60]*tmp[162]+tmp[61]*tmp[161]+tmp[62]*tmp[160]+tmp[63]*tmp[159]+tmp[64]*tmp[158]+tmp[65]*tmp[157]+tmp[66]*tmp[156]+tmp[67]*tmp[155]+tmp[68]*tmp[154]+tmp[69]*tmp[153]+tmp[70]*tmp[152]+tmp[71]*tmp[151]+tmp[72]*tmp[150]+tmp[73]*tmp[149]+tmp[74]*tmp[148]+tmp[75]*tmp[147]+tmp[76]*tmp[146]+tmp[77]*tmp[145]+tmp[78]*tmp[144]+tmp[79]*tmp[143]+tmp[80]*tmp[142]+tmp[81]*tmp[141]+tmp[82]*tmp[140]+tmp[83]*tmp[139]+tmp[84]*tmp[138]+tmp[85]*tmp[137]+tmp[86]*tmp[136]+tmp[87]*tmp[135]+tmp[88]*tmp[134]+tmp[89]*tmp[133]+tmp[90]*tmp[132]+tmp[91]*tmp[131]+tmp[92]*tmp[130]+tmp[93]*tmp[129]+tmp[94]*tmp[128]+tmp[95]*tmp[127]+tmp[96]*tmp[126]+tmp[97]*tmp[125]+tmp[98]*tmp[124]+tmp[99]*tmp[123];
				ans[123]<=tmp[24]*tmp[199]+tmp[25]*tmp[198]+tmp[26]*tmp[197]+tmp[27]*tmp[196]+tmp[28]*tmp[195]+tmp[29]*tmp[194]+tmp[30]*tmp[193]+tmp[31]*tmp[192]+tmp[32]*tmp[191]+tmp[33]*tmp[190]+tmp[34]*tmp[189]+tmp[35]*tmp[188]+tmp[36]*tmp[187]+tmp[37]*tmp[186]+tmp[38]*tmp[185]+tmp[39]*tmp[184]+tmp[40]*tmp[183]+tmp[41]*tmp[182]+tmp[42]*tmp[181]+tmp[43]*tmp[180]+tmp[44]*tmp[179]+tmp[45]*tmp[178]+tmp[46]*tmp[177]+tmp[47]*tmp[176]+tmp[48]*tmp[175]+tmp[49]*tmp[174]+tmp[50]*tmp[173]+tmp[51]*tmp[172]+tmp[52]*tmp[171]+tmp[53]*tmp[170]+tmp[54]*tmp[169]+tmp[55]*tmp[168]+tmp[56]*tmp[167]+tmp[57]*tmp[166]+tmp[58]*tmp[165]+tmp[59]*tmp[164]+tmp[60]*tmp[163]+tmp[61]*tmp[162]+tmp[62]*tmp[161]+tmp[63]*tmp[160]+tmp[64]*tmp[159]+tmp[65]*tmp[158]+tmp[66]*tmp[157]+tmp[67]*tmp[156]+tmp[68]*tmp[155]+tmp[69]*tmp[154]+tmp[70]*tmp[153]+tmp[71]*tmp[152]+tmp[72]*tmp[151]+tmp[73]*tmp[150]+tmp[74]*tmp[149]+tmp[75]*tmp[148]+tmp[76]*tmp[147]+tmp[77]*tmp[146]+tmp[78]*tmp[145]+tmp[79]*tmp[144]+tmp[80]*tmp[143]+tmp[81]*tmp[142]+tmp[82]*tmp[141]+tmp[83]*tmp[140]+tmp[84]*tmp[139]+tmp[85]*tmp[138]+tmp[86]*tmp[137]+tmp[87]*tmp[136]+tmp[88]*tmp[135]+tmp[89]*tmp[134]+tmp[90]*tmp[133]+tmp[91]*tmp[132]+tmp[92]*tmp[131]+tmp[93]*tmp[130]+tmp[94]*tmp[129]+tmp[95]*tmp[128]+tmp[96]*tmp[127]+tmp[97]*tmp[126]+tmp[98]*tmp[125]+tmp[99]*tmp[124];
				ans[124]<=tmp[25]*tmp[199]+tmp[26]*tmp[198]+tmp[27]*tmp[197]+tmp[28]*tmp[196]+tmp[29]*tmp[195]+tmp[30]*tmp[194]+tmp[31]*tmp[193]+tmp[32]*tmp[192]+tmp[33]*tmp[191]+tmp[34]*tmp[190]+tmp[35]*tmp[189]+tmp[36]*tmp[188]+tmp[37]*tmp[187]+tmp[38]*tmp[186]+tmp[39]*tmp[185]+tmp[40]*tmp[184]+tmp[41]*tmp[183]+tmp[42]*tmp[182]+tmp[43]*tmp[181]+tmp[44]*tmp[180]+tmp[45]*tmp[179]+tmp[46]*tmp[178]+tmp[47]*tmp[177]+tmp[48]*tmp[176]+tmp[49]*tmp[175]+tmp[50]*tmp[174]+tmp[51]*tmp[173]+tmp[52]*tmp[172]+tmp[53]*tmp[171]+tmp[54]*tmp[170]+tmp[55]*tmp[169]+tmp[56]*tmp[168]+tmp[57]*tmp[167]+tmp[58]*tmp[166]+tmp[59]*tmp[165]+tmp[60]*tmp[164]+tmp[61]*tmp[163]+tmp[62]*tmp[162]+tmp[63]*tmp[161]+tmp[64]*tmp[160]+tmp[65]*tmp[159]+tmp[66]*tmp[158]+tmp[67]*tmp[157]+tmp[68]*tmp[156]+tmp[69]*tmp[155]+tmp[70]*tmp[154]+tmp[71]*tmp[153]+tmp[72]*tmp[152]+tmp[73]*tmp[151]+tmp[74]*tmp[150]+tmp[75]*tmp[149]+tmp[76]*tmp[148]+tmp[77]*tmp[147]+tmp[78]*tmp[146]+tmp[79]*tmp[145]+tmp[80]*tmp[144]+tmp[81]*tmp[143]+tmp[82]*tmp[142]+tmp[83]*tmp[141]+tmp[84]*tmp[140]+tmp[85]*tmp[139]+tmp[86]*tmp[138]+tmp[87]*tmp[137]+tmp[88]*tmp[136]+tmp[89]*tmp[135]+tmp[90]*tmp[134]+tmp[91]*tmp[133]+tmp[92]*tmp[132]+tmp[93]*tmp[131]+tmp[94]*tmp[130]+tmp[95]*tmp[129]+tmp[96]*tmp[128]+tmp[97]*tmp[127]+tmp[98]*tmp[126]+tmp[99]*tmp[125];
				ans[125]<=tmp[26]*tmp[199]+tmp[27]*tmp[198]+tmp[28]*tmp[197]+tmp[29]*tmp[196]+tmp[30]*tmp[195]+tmp[31]*tmp[194]+tmp[32]*tmp[193]+tmp[33]*tmp[192]+tmp[34]*tmp[191]+tmp[35]*tmp[190]+tmp[36]*tmp[189]+tmp[37]*tmp[188]+tmp[38]*tmp[187]+tmp[39]*tmp[186]+tmp[40]*tmp[185]+tmp[41]*tmp[184]+tmp[42]*tmp[183]+tmp[43]*tmp[182]+tmp[44]*tmp[181]+tmp[45]*tmp[180]+tmp[46]*tmp[179]+tmp[47]*tmp[178]+tmp[48]*tmp[177]+tmp[49]*tmp[176]+tmp[50]*tmp[175]+tmp[51]*tmp[174]+tmp[52]*tmp[173]+tmp[53]*tmp[172]+tmp[54]*tmp[171]+tmp[55]*tmp[170]+tmp[56]*tmp[169]+tmp[57]*tmp[168]+tmp[58]*tmp[167]+tmp[59]*tmp[166]+tmp[60]*tmp[165]+tmp[61]*tmp[164]+tmp[62]*tmp[163]+tmp[63]*tmp[162]+tmp[64]*tmp[161]+tmp[65]*tmp[160]+tmp[66]*tmp[159]+tmp[67]*tmp[158]+tmp[68]*tmp[157]+tmp[69]*tmp[156]+tmp[70]*tmp[155]+tmp[71]*tmp[154]+tmp[72]*tmp[153]+tmp[73]*tmp[152]+tmp[74]*tmp[151]+tmp[75]*tmp[150]+tmp[76]*tmp[149]+tmp[77]*tmp[148]+tmp[78]*tmp[147]+tmp[79]*tmp[146]+tmp[80]*tmp[145]+tmp[81]*tmp[144]+tmp[82]*tmp[143]+tmp[83]*tmp[142]+tmp[84]*tmp[141]+tmp[85]*tmp[140]+tmp[86]*tmp[139]+tmp[87]*tmp[138]+tmp[88]*tmp[137]+tmp[89]*tmp[136]+tmp[90]*tmp[135]+tmp[91]*tmp[134]+tmp[92]*tmp[133]+tmp[93]*tmp[132]+tmp[94]*tmp[131]+tmp[95]*tmp[130]+tmp[96]*tmp[129]+tmp[97]*tmp[128]+tmp[98]*tmp[127]+tmp[99]*tmp[126];
				ans[126]<=tmp[27]*tmp[199]+tmp[28]*tmp[198]+tmp[29]*tmp[197]+tmp[30]*tmp[196]+tmp[31]*tmp[195]+tmp[32]*tmp[194]+tmp[33]*tmp[193]+tmp[34]*tmp[192]+tmp[35]*tmp[191]+tmp[36]*tmp[190]+tmp[37]*tmp[189]+tmp[38]*tmp[188]+tmp[39]*tmp[187]+tmp[40]*tmp[186]+tmp[41]*tmp[185]+tmp[42]*tmp[184]+tmp[43]*tmp[183]+tmp[44]*tmp[182]+tmp[45]*tmp[181]+tmp[46]*tmp[180]+tmp[47]*tmp[179]+tmp[48]*tmp[178]+tmp[49]*tmp[177]+tmp[50]*tmp[176]+tmp[51]*tmp[175]+tmp[52]*tmp[174]+tmp[53]*tmp[173]+tmp[54]*tmp[172]+tmp[55]*tmp[171]+tmp[56]*tmp[170]+tmp[57]*tmp[169]+tmp[58]*tmp[168]+tmp[59]*tmp[167]+tmp[60]*tmp[166]+tmp[61]*tmp[165]+tmp[62]*tmp[164]+tmp[63]*tmp[163]+tmp[64]*tmp[162]+tmp[65]*tmp[161]+tmp[66]*tmp[160]+tmp[67]*tmp[159]+tmp[68]*tmp[158]+tmp[69]*tmp[157]+tmp[70]*tmp[156]+tmp[71]*tmp[155]+tmp[72]*tmp[154]+tmp[73]*tmp[153]+tmp[74]*tmp[152]+tmp[75]*tmp[151]+tmp[76]*tmp[150]+tmp[77]*tmp[149]+tmp[78]*tmp[148]+tmp[79]*tmp[147]+tmp[80]*tmp[146]+tmp[81]*tmp[145]+tmp[82]*tmp[144]+tmp[83]*tmp[143]+tmp[84]*tmp[142]+tmp[85]*tmp[141]+tmp[86]*tmp[140]+tmp[87]*tmp[139]+tmp[88]*tmp[138]+tmp[89]*tmp[137]+tmp[90]*tmp[136]+tmp[91]*tmp[135]+tmp[92]*tmp[134]+tmp[93]*tmp[133]+tmp[94]*tmp[132]+tmp[95]*tmp[131]+tmp[96]*tmp[130]+tmp[97]*tmp[129]+tmp[98]*tmp[128]+tmp[99]*tmp[127];
				ans[127]<=tmp[28]*tmp[199]+tmp[29]*tmp[198]+tmp[30]*tmp[197]+tmp[31]*tmp[196]+tmp[32]*tmp[195]+tmp[33]*tmp[194]+tmp[34]*tmp[193]+tmp[35]*tmp[192]+tmp[36]*tmp[191]+tmp[37]*tmp[190]+tmp[38]*tmp[189]+tmp[39]*tmp[188]+tmp[40]*tmp[187]+tmp[41]*tmp[186]+tmp[42]*tmp[185]+tmp[43]*tmp[184]+tmp[44]*tmp[183]+tmp[45]*tmp[182]+tmp[46]*tmp[181]+tmp[47]*tmp[180]+tmp[48]*tmp[179]+tmp[49]*tmp[178]+tmp[50]*tmp[177]+tmp[51]*tmp[176]+tmp[52]*tmp[175]+tmp[53]*tmp[174]+tmp[54]*tmp[173]+tmp[55]*tmp[172]+tmp[56]*tmp[171]+tmp[57]*tmp[170]+tmp[58]*tmp[169]+tmp[59]*tmp[168]+tmp[60]*tmp[167]+tmp[61]*tmp[166]+tmp[62]*tmp[165]+tmp[63]*tmp[164]+tmp[64]*tmp[163]+tmp[65]*tmp[162]+tmp[66]*tmp[161]+tmp[67]*tmp[160]+tmp[68]*tmp[159]+tmp[69]*tmp[158]+tmp[70]*tmp[157]+tmp[71]*tmp[156]+tmp[72]*tmp[155]+tmp[73]*tmp[154]+tmp[74]*tmp[153]+tmp[75]*tmp[152]+tmp[76]*tmp[151]+tmp[77]*tmp[150]+tmp[78]*tmp[149]+tmp[79]*tmp[148]+tmp[80]*tmp[147]+tmp[81]*tmp[146]+tmp[82]*tmp[145]+tmp[83]*tmp[144]+tmp[84]*tmp[143]+tmp[85]*tmp[142]+tmp[86]*tmp[141]+tmp[87]*tmp[140]+tmp[88]*tmp[139]+tmp[89]*tmp[138]+tmp[90]*tmp[137]+tmp[91]*tmp[136]+tmp[92]*tmp[135]+tmp[93]*tmp[134]+tmp[94]*tmp[133]+tmp[95]*tmp[132]+tmp[96]*tmp[131]+tmp[97]*tmp[130]+tmp[98]*tmp[129]+tmp[99]*tmp[128];
				ans[128]<=tmp[29]*tmp[199]+tmp[30]*tmp[198]+tmp[31]*tmp[197]+tmp[32]*tmp[196]+tmp[33]*tmp[195]+tmp[34]*tmp[194]+tmp[35]*tmp[193]+tmp[36]*tmp[192]+tmp[37]*tmp[191]+tmp[38]*tmp[190]+tmp[39]*tmp[189]+tmp[40]*tmp[188]+tmp[41]*tmp[187]+tmp[42]*tmp[186]+tmp[43]*tmp[185]+tmp[44]*tmp[184]+tmp[45]*tmp[183]+tmp[46]*tmp[182]+tmp[47]*tmp[181]+tmp[48]*tmp[180]+tmp[49]*tmp[179]+tmp[50]*tmp[178]+tmp[51]*tmp[177]+tmp[52]*tmp[176]+tmp[53]*tmp[175]+tmp[54]*tmp[174]+tmp[55]*tmp[173]+tmp[56]*tmp[172]+tmp[57]*tmp[171]+tmp[58]*tmp[170]+tmp[59]*tmp[169]+tmp[60]*tmp[168]+tmp[61]*tmp[167]+tmp[62]*tmp[166]+tmp[63]*tmp[165]+tmp[64]*tmp[164]+tmp[65]*tmp[163]+tmp[66]*tmp[162]+tmp[67]*tmp[161]+tmp[68]*tmp[160]+tmp[69]*tmp[159]+tmp[70]*tmp[158]+tmp[71]*tmp[157]+tmp[72]*tmp[156]+tmp[73]*tmp[155]+tmp[74]*tmp[154]+tmp[75]*tmp[153]+tmp[76]*tmp[152]+tmp[77]*tmp[151]+tmp[78]*tmp[150]+tmp[79]*tmp[149]+tmp[80]*tmp[148]+tmp[81]*tmp[147]+tmp[82]*tmp[146]+tmp[83]*tmp[145]+tmp[84]*tmp[144]+tmp[85]*tmp[143]+tmp[86]*tmp[142]+tmp[87]*tmp[141]+tmp[88]*tmp[140]+tmp[89]*tmp[139]+tmp[90]*tmp[138]+tmp[91]*tmp[137]+tmp[92]*tmp[136]+tmp[93]*tmp[135]+tmp[94]*tmp[134]+tmp[95]*tmp[133]+tmp[96]*tmp[132]+tmp[97]*tmp[131]+tmp[98]*tmp[130]+tmp[99]*tmp[129];
				ans[129]<=tmp[30]*tmp[199]+tmp[31]*tmp[198]+tmp[32]*tmp[197]+tmp[33]*tmp[196]+tmp[34]*tmp[195]+tmp[35]*tmp[194]+tmp[36]*tmp[193]+tmp[37]*tmp[192]+tmp[38]*tmp[191]+tmp[39]*tmp[190]+tmp[40]*tmp[189]+tmp[41]*tmp[188]+tmp[42]*tmp[187]+tmp[43]*tmp[186]+tmp[44]*tmp[185]+tmp[45]*tmp[184]+tmp[46]*tmp[183]+tmp[47]*tmp[182]+tmp[48]*tmp[181]+tmp[49]*tmp[180]+tmp[50]*tmp[179]+tmp[51]*tmp[178]+tmp[52]*tmp[177]+tmp[53]*tmp[176]+tmp[54]*tmp[175]+tmp[55]*tmp[174]+tmp[56]*tmp[173]+tmp[57]*tmp[172]+tmp[58]*tmp[171]+tmp[59]*tmp[170]+tmp[60]*tmp[169]+tmp[61]*tmp[168]+tmp[62]*tmp[167]+tmp[63]*tmp[166]+tmp[64]*tmp[165]+tmp[65]*tmp[164]+tmp[66]*tmp[163]+tmp[67]*tmp[162]+tmp[68]*tmp[161]+tmp[69]*tmp[160]+tmp[70]*tmp[159]+tmp[71]*tmp[158]+tmp[72]*tmp[157]+tmp[73]*tmp[156]+tmp[74]*tmp[155]+tmp[75]*tmp[154]+tmp[76]*tmp[153]+tmp[77]*tmp[152]+tmp[78]*tmp[151]+tmp[79]*tmp[150]+tmp[80]*tmp[149]+tmp[81]*tmp[148]+tmp[82]*tmp[147]+tmp[83]*tmp[146]+tmp[84]*tmp[145]+tmp[85]*tmp[144]+tmp[86]*tmp[143]+tmp[87]*tmp[142]+tmp[88]*tmp[141]+tmp[89]*tmp[140]+tmp[90]*tmp[139]+tmp[91]*tmp[138]+tmp[92]*tmp[137]+tmp[93]*tmp[136]+tmp[94]*tmp[135]+tmp[95]*tmp[134]+tmp[96]*tmp[133]+tmp[97]*tmp[132]+tmp[98]*tmp[131]+tmp[99]*tmp[130];
				ans[130]<=tmp[31]*tmp[199]+tmp[32]*tmp[198]+tmp[33]*tmp[197]+tmp[34]*tmp[196]+tmp[35]*tmp[195]+tmp[36]*tmp[194]+tmp[37]*tmp[193]+tmp[38]*tmp[192]+tmp[39]*tmp[191]+tmp[40]*tmp[190]+tmp[41]*tmp[189]+tmp[42]*tmp[188]+tmp[43]*tmp[187]+tmp[44]*tmp[186]+tmp[45]*tmp[185]+tmp[46]*tmp[184]+tmp[47]*tmp[183]+tmp[48]*tmp[182]+tmp[49]*tmp[181]+tmp[50]*tmp[180]+tmp[51]*tmp[179]+tmp[52]*tmp[178]+tmp[53]*tmp[177]+tmp[54]*tmp[176]+tmp[55]*tmp[175]+tmp[56]*tmp[174]+tmp[57]*tmp[173]+tmp[58]*tmp[172]+tmp[59]*tmp[171]+tmp[60]*tmp[170]+tmp[61]*tmp[169]+tmp[62]*tmp[168]+tmp[63]*tmp[167]+tmp[64]*tmp[166]+tmp[65]*tmp[165]+tmp[66]*tmp[164]+tmp[67]*tmp[163]+tmp[68]*tmp[162]+tmp[69]*tmp[161]+tmp[70]*tmp[160]+tmp[71]*tmp[159]+tmp[72]*tmp[158]+tmp[73]*tmp[157]+tmp[74]*tmp[156]+tmp[75]*tmp[155]+tmp[76]*tmp[154]+tmp[77]*tmp[153]+tmp[78]*tmp[152]+tmp[79]*tmp[151]+tmp[80]*tmp[150]+tmp[81]*tmp[149]+tmp[82]*tmp[148]+tmp[83]*tmp[147]+tmp[84]*tmp[146]+tmp[85]*tmp[145]+tmp[86]*tmp[144]+tmp[87]*tmp[143]+tmp[88]*tmp[142]+tmp[89]*tmp[141]+tmp[90]*tmp[140]+tmp[91]*tmp[139]+tmp[92]*tmp[138]+tmp[93]*tmp[137]+tmp[94]*tmp[136]+tmp[95]*tmp[135]+tmp[96]*tmp[134]+tmp[97]*tmp[133]+tmp[98]*tmp[132]+tmp[99]*tmp[131];
				ans[131]<=tmp[32]*tmp[199]+tmp[33]*tmp[198]+tmp[34]*tmp[197]+tmp[35]*tmp[196]+tmp[36]*tmp[195]+tmp[37]*tmp[194]+tmp[38]*tmp[193]+tmp[39]*tmp[192]+tmp[40]*tmp[191]+tmp[41]*tmp[190]+tmp[42]*tmp[189]+tmp[43]*tmp[188]+tmp[44]*tmp[187]+tmp[45]*tmp[186]+tmp[46]*tmp[185]+tmp[47]*tmp[184]+tmp[48]*tmp[183]+tmp[49]*tmp[182]+tmp[50]*tmp[181]+tmp[51]*tmp[180]+tmp[52]*tmp[179]+tmp[53]*tmp[178]+tmp[54]*tmp[177]+tmp[55]*tmp[176]+tmp[56]*tmp[175]+tmp[57]*tmp[174]+tmp[58]*tmp[173]+tmp[59]*tmp[172]+tmp[60]*tmp[171]+tmp[61]*tmp[170]+tmp[62]*tmp[169]+tmp[63]*tmp[168]+tmp[64]*tmp[167]+tmp[65]*tmp[166]+tmp[66]*tmp[165]+tmp[67]*tmp[164]+tmp[68]*tmp[163]+tmp[69]*tmp[162]+tmp[70]*tmp[161]+tmp[71]*tmp[160]+tmp[72]*tmp[159]+tmp[73]*tmp[158]+tmp[74]*tmp[157]+tmp[75]*tmp[156]+tmp[76]*tmp[155]+tmp[77]*tmp[154]+tmp[78]*tmp[153]+tmp[79]*tmp[152]+tmp[80]*tmp[151]+tmp[81]*tmp[150]+tmp[82]*tmp[149]+tmp[83]*tmp[148]+tmp[84]*tmp[147]+tmp[85]*tmp[146]+tmp[86]*tmp[145]+tmp[87]*tmp[144]+tmp[88]*tmp[143]+tmp[89]*tmp[142]+tmp[90]*tmp[141]+tmp[91]*tmp[140]+tmp[92]*tmp[139]+tmp[93]*tmp[138]+tmp[94]*tmp[137]+tmp[95]*tmp[136]+tmp[96]*tmp[135]+tmp[97]*tmp[134]+tmp[98]*tmp[133]+tmp[99]*tmp[132];
				ans[132]<=tmp[33]*tmp[199]+tmp[34]*tmp[198]+tmp[35]*tmp[197]+tmp[36]*tmp[196]+tmp[37]*tmp[195]+tmp[38]*tmp[194]+tmp[39]*tmp[193]+tmp[40]*tmp[192]+tmp[41]*tmp[191]+tmp[42]*tmp[190]+tmp[43]*tmp[189]+tmp[44]*tmp[188]+tmp[45]*tmp[187]+tmp[46]*tmp[186]+tmp[47]*tmp[185]+tmp[48]*tmp[184]+tmp[49]*tmp[183]+tmp[50]*tmp[182]+tmp[51]*tmp[181]+tmp[52]*tmp[180]+tmp[53]*tmp[179]+tmp[54]*tmp[178]+tmp[55]*tmp[177]+tmp[56]*tmp[176]+tmp[57]*tmp[175]+tmp[58]*tmp[174]+tmp[59]*tmp[173]+tmp[60]*tmp[172]+tmp[61]*tmp[171]+tmp[62]*tmp[170]+tmp[63]*tmp[169]+tmp[64]*tmp[168]+tmp[65]*tmp[167]+tmp[66]*tmp[166]+tmp[67]*tmp[165]+tmp[68]*tmp[164]+tmp[69]*tmp[163]+tmp[70]*tmp[162]+tmp[71]*tmp[161]+tmp[72]*tmp[160]+tmp[73]*tmp[159]+tmp[74]*tmp[158]+tmp[75]*tmp[157]+tmp[76]*tmp[156]+tmp[77]*tmp[155]+tmp[78]*tmp[154]+tmp[79]*tmp[153]+tmp[80]*tmp[152]+tmp[81]*tmp[151]+tmp[82]*tmp[150]+tmp[83]*tmp[149]+tmp[84]*tmp[148]+tmp[85]*tmp[147]+tmp[86]*tmp[146]+tmp[87]*tmp[145]+tmp[88]*tmp[144]+tmp[89]*tmp[143]+tmp[90]*tmp[142]+tmp[91]*tmp[141]+tmp[92]*tmp[140]+tmp[93]*tmp[139]+tmp[94]*tmp[138]+tmp[95]*tmp[137]+tmp[96]*tmp[136]+tmp[97]*tmp[135]+tmp[98]*tmp[134]+tmp[99]*tmp[133];
				ans[133]<=tmp[34]*tmp[199]+tmp[35]*tmp[198]+tmp[36]*tmp[197]+tmp[37]*tmp[196]+tmp[38]*tmp[195]+tmp[39]*tmp[194]+tmp[40]*tmp[193]+tmp[41]*tmp[192]+tmp[42]*tmp[191]+tmp[43]*tmp[190]+tmp[44]*tmp[189]+tmp[45]*tmp[188]+tmp[46]*tmp[187]+tmp[47]*tmp[186]+tmp[48]*tmp[185]+tmp[49]*tmp[184]+tmp[50]*tmp[183]+tmp[51]*tmp[182]+tmp[52]*tmp[181]+tmp[53]*tmp[180]+tmp[54]*tmp[179]+tmp[55]*tmp[178]+tmp[56]*tmp[177]+tmp[57]*tmp[176]+tmp[58]*tmp[175]+tmp[59]*tmp[174]+tmp[60]*tmp[173]+tmp[61]*tmp[172]+tmp[62]*tmp[171]+tmp[63]*tmp[170]+tmp[64]*tmp[169]+tmp[65]*tmp[168]+tmp[66]*tmp[167]+tmp[67]*tmp[166]+tmp[68]*tmp[165]+tmp[69]*tmp[164]+tmp[70]*tmp[163]+tmp[71]*tmp[162]+tmp[72]*tmp[161]+tmp[73]*tmp[160]+tmp[74]*tmp[159]+tmp[75]*tmp[158]+tmp[76]*tmp[157]+tmp[77]*tmp[156]+tmp[78]*tmp[155]+tmp[79]*tmp[154]+tmp[80]*tmp[153]+tmp[81]*tmp[152]+tmp[82]*tmp[151]+tmp[83]*tmp[150]+tmp[84]*tmp[149]+tmp[85]*tmp[148]+tmp[86]*tmp[147]+tmp[87]*tmp[146]+tmp[88]*tmp[145]+tmp[89]*tmp[144]+tmp[90]*tmp[143]+tmp[91]*tmp[142]+tmp[92]*tmp[141]+tmp[93]*tmp[140]+tmp[94]*tmp[139]+tmp[95]*tmp[138]+tmp[96]*tmp[137]+tmp[97]*tmp[136]+tmp[98]*tmp[135]+tmp[99]*tmp[134];
				ans[134]<=tmp[35]*tmp[199]+tmp[36]*tmp[198]+tmp[37]*tmp[197]+tmp[38]*tmp[196]+tmp[39]*tmp[195]+tmp[40]*tmp[194]+tmp[41]*tmp[193]+tmp[42]*tmp[192]+tmp[43]*tmp[191]+tmp[44]*tmp[190]+tmp[45]*tmp[189]+tmp[46]*tmp[188]+tmp[47]*tmp[187]+tmp[48]*tmp[186]+tmp[49]*tmp[185]+tmp[50]*tmp[184]+tmp[51]*tmp[183]+tmp[52]*tmp[182]+tmp[53]*tmp[181]+tmp[54]*tmp[180]+tmp[55]*tmp[179]+tmp[56]*tmp[178]+tmp[57]*tmp[177]+tmp[58]*tmp[176]+tmp[59]*tmp[175]+tmp[60]*tmp[174]+tmp[61]*tmp[173]+tmp[62]*tmp[172]+tmp[63]*tmp[171]+tmp[64]*tmp[170]+tmp[65]*tmp[169]+tmp[66]*tmp[168]+tmp[67]*tmp[167]+tmp[68]*tmp[166]+tmp[69]*tmp[165]+tmp[70]*tmp[164]+tmp[71]*tmp[163]+tmp[72]*tmp[162]+tmp[73]*tmp[161]+tmp[74]*tmp[160]+tmp[75]*tmp[159]+tmp[76]*tmp[158]+tmp[77]*tmp[157]+tmp[78]*tmp[156]+tmp[79]*tmp[155]+tmp[80]*tmp[154]+tmp[81]*tmp[153]+tmp[82]*tmp[152]+tmp[83]*tmp[151]+tmp[84]*tmp[150]+tmp[85]*tmp[149]+tmp[86]*tmp[148]+tmp[87]*tmp[147]+tmp[88]*tmp[146]+tmp[89]*tmp[145]+tmp[90]*tmp[144]+tmp[91]*tmp[143]+tmp[92]*tmp[142]+tmp[93]*tmp[141]+tmp[94]*tmp[140]+tmp[95]*tmp[139]+tmp[96]*tmp[138]+tmp[97]*tmp[137]+tmp[98]*tmp[136]+tmp[99]*tmp[135];
				ans[135]<=tmp[36]*tmp[199]+tmp[37]*tmp[198]+tmp[38]*tmp[197]+tmp[39]*tmp[196]+tmp[40]*tmp[195]+tmp[41]*tmp[194]+tmp[42]*tmp[193]+tmp[43]*tmp[192]+tmp[44]*tmp[191]+tmp[45]*tmp[190]+tmp[46]*tmp[189]+tmp[47]*tmp[188]+tmp[48]*tmp[187]+tmp[49]*tmp[186]+tmp[50]*tmp[185]+tmp[51]*tmp[184]+tmp[52]*tmp[183]+tmp[53]*tmp[182]+tmp[54]*tmp[181]+tmp[55]*tmp[180]+tmp[56]*tmp[179]+tmp[57]*tmp[178]+tmp[58]*tmp[177]+tmp[59]*tmp[176]+tmp[60]*tmp[175]+tmp[61]*tmp[174]+tmp[62]*tmp[173]+tmp[63]*tmp[172]+tmp[64]*tmp[171]+tmp[65]*tmp[170]+tmp[66]*tmp[169]+tmp[67]*tmp[168]+tmp[68]*tmp[167]+tmp[69]*tmp[166]+tmp[70]*tmp[165]+tmp[71]*tmp[164]+tmp[72]*tmp[163]+tmp[73]*tmp[162]+tmp[74]*tmp[161]+tmp[75]*tmp[160]+tmp[76]*tmp[159]+tmp[77]*tmp[158]+tmp[78]*tmp[157]+tmp[79]*tmp[156]+tmp[80]*tmp[155]+tmp[81]*tmp[154]+tmp[82]*tmp[153]+tmp[83]*tmp[152]+tmp[84]*tmp[151]+tmp[85]*tmp[150]+tmp[86]*tmp[149]+tmp[87]*tmp[148]+tmp[88]*tmp[147]+tmp[89]*tmp[146]+tmp[90]*tmp[145]+tmp[91]*tmp[144]+tmp[92]*tmp[143]+tmp[93]*tmp[142]+tmp[94]*tmp[141]+tmp[95]*tmp[140]+tmp[96]*tmp[139]+tmp[97]*tmp[138]+tmp[98]*tmp[137]+tmp[99]*tmp[136];
				ans[136]<=tmp[37]*tmp[199]+tmp[38]*tmp[198]+tmp[39]*tmp[197]+tmp[40]*tmp[196]+tmp[41]*tmp[195]+tmp[42]*tmp[194]+tmp[43]*tmp[193]+tmp[44]*tmp[192]+tmp[45]*tmp[191]+tmp[46]*tmp[190]+tmp[47]*tmp[189]+tmp[48]*tmp[188]+tmp[49]*tmp[187]+tmp[50]*tmp[186]+tmp[51]*tmp[185]+tmp[52]*tmp[184]+tmp[53]*tmp[183]+tmp[54]*tmp[182]+tmp[55]*tmp[181]+tmp[56]*tmp[180]+tmp[57]*tmp[179]+tmp[58]*tmp[178]+tmp[59]*tmp[177]+tmp[60]*tmp[176]+tmp[61]*tmp[175]+tmp[62]*tmp[174]+tmp[63]*tmp[173]+tmp[64]*tmp[172]+tmp[65]*tmp[171]+tmp[66]*tmp[170]+tmp[67]*tmp[169]+tmp[68]*tmp[168]+tmp[69]*tmp[167]+tmp[70]*tmp[166]+tmp[71]*tmp[165]+tmp[72]*tmp[164]+tmp[73]*tmp[163]+tmp[74]*tmp[162]+tmp[75]*tmp[161]+tmp[76]*tmp[160]+tmp[77]*tmp[159]+tmp[78]*tmp[158]+tmp[79]*tmp[157]+tmp[80]*tmp[156]+tmp[81]*tmp[155]+tmp[82]*tmp[154]+tmp[83]*tmp[153]+tmp[84]*tmp[152]+tmp[85]*tmp[151]+tmp[86]*tmp[150]+tmp[87]*tmp[149]+tmp[88]*tmp[148]+tmp[89]*tmp[147]+tmp[90]*tmp[146]+tmp[91]*tmp[145]+tmp[92]*tmp[144]+tmp[93]*tmp[143]+tmp[94]*tmp[142]+tmp[95]*tmp[141]+tmp[96]*tmp[140]+tmp[97]*tmp[139]+tmp[98]*tmp[138]+tmp[99]*tmp[137];
				ans[137]<=tmp[38]*tmp[199]+tmp[39]*tmp[198]+tmp[40]*tmp[197]+tmp[41]*tmp[196]+tmp[42]*tmp[195]+tmp[43]*tmp[194]+tmp[44]*tmp[193]+tmp[45]*tmp[192]+tmp[46]*tmp[191]+tmp[47]*tmp[190]+tmp[48]*tmp[189]+tmp[49]*tmp[188]+tmp[50]*tmp[187]+tmp[51]*tmp[186]+tmp[52]*tmp[185]+tmp[53]*tmp[184]+tmp[54]*tmp[183]+tmp[55]*tmp[182]+tmp[56]*tmp[181]+tmp[57]*tmp[180]+tmp[58]*tmp[179]+tmp[59]*tmp[178]+tmp[60]*tmp[177]+tmp[61]*tmp[176]+tmp[62]*tmp[175]+tmp[63]*tmp[174]+tmp[64]*tmp[173]+tmp[65]*tmp[172]+tmp[66]*tmp[171]+tmp[67]*tmp[170]+tmp[68]*tmp[169]+tmp[69]*tmp[168]+tmp[70]*tmp[167]+tmp[71]*tmp[166]+tmp[72]*tmp[165]+tmp[73]*tmp[164]+tmp[74]*tmp[163]+tmp[75]*tmp[162]+tmp[76]*tmp[161]+tmp[77]*tmp[160]+tmp[78]*tmp[159]+tmp[79]*tmp[158]+tmp[80]*tmp[157]+tmp[81]*tmp[156]+tmp[82]*tmp[155]+tmp[83]*tmp[154]+tmp[84]*tmp[153]+tmp[85]*tmp[152]+tmp[86]*tmp[151]+tmp[87]*tmp[150]+tmp[88]*tmp[149]+tmp[89]*tmp[148]+tmp[90]*tmp[147]+tmp[91]*tmp[146]+tmp[92]*tmp[145]+tmp[93]*tmp[144]+tmp[94]*tmp[143]+tmp[95]*tmp[142]+tmp[96]*tmp[141]+tmp[97]*tmp[140]+tmp[98]*tmp[139]+tmp[99]*tmp[138];
				ans[138]<=tmp[39]*tmp[199]+tmp[40]*tmp[198]+tmp[41]*tmp[197]+tmp[42]*tmp[196]+tmp[43]*tmp[195]+tmp[44]*tmp[194]+tmp[45]*tmp[193]+tmp[46]*tmp[192]+tmp[47]*tmp[191]+tmp[48]*tmp[190]+tmp[49]*tmp[189]+tmp[50]*tmp[188]+tmp[51]*tmp[187]+tmp[52]*tmp[186]+tmp[53]*tmp[185]+tmp[54]*tmp[184]+tmp[55]*tmp[183]+tmp[56]*tmp[182]+tmp[57]*tmp[181]+tmp[58]*tmp[180]+tmp[59]*tmp[179]+tmp[60]*tmp[178]+tmp[61]*tmp[177]+tmp[62]*tmp[176]+tmp[63]*tmp[175]+tmp[64]*tmp[174]+tmp[65]*tmp[173]+tmp[66]*tmp[172]+tmp[67]*tmp[171]+tmp[68]*tmp[170]+tmp[69]*tmp[169]+tmp[70]*tmp[168]+tmp[71]*tmp[167]+tmp[72]*tmp[166]+tmp[73]*tmp[165]+tmp[74]*tmp[164]+tmp[75]*tmp[163]+tmp[76]*tmp[162]+tmp[77]*tmp[161]+tmp[78]*tmp[160]+tmp[79]*tmp[159]+tmp[80]*tmp[158]+tmp[81]*tmp[157]+tmp[82]*tmp[156]+tmp[83]*tmp[155]+tmp[84]*tmp[154]+tmp[85]*tmp[153]+tmp[86]*tmp[152]+tmp[87]*tmp[151]+tmp[88]*tmp[150]+tmp[89]*tmp[149]+tmp[90]*tmp[148]+tmp[91]*tmp[147]+tmp[92]*tmp[146]+tmp[93]*tmp[145]+tmp[94]*tmp[144]+tmp[95]*tmp[143]+tmp[96]*tmp[142]+tmp[97]*tmp[141]+tmp[98]*tmp[140]+tmp[99]*tmp[139];
				ans[139]<=tmp[40]*tmp[199]+tmp[41]*tmp[198]+tmp[42]*tmp[197]+tmp[43]*tmp[196]+tmp[44]*tmp[195]+tmp[45]*tmp[194]+tmp[46]*tmp[193]+tmp[47]*tmp[192]+tmp[48]*tmp[191]+tmp[49]*tmp[190]+tmp[50]*tmp[189]+tmp[51]*tmp[188]+tmp[52]*tmp[187]+tmp[53]*tmp[186]+tmp[54]*tmp[185]+tmp[55]*tmp[184]+tmp[56]*tmp[183]+tmp[57]*tmp[182]+tmp[58]*tmp[181]+tmp[59]*tmp[180]+tmp[60]*tmp[179]+tmp[61]*tmp[178]+tmp[62]*tmp[177]+tmp[63]*tmp[176]+tmp[64]*tmp[175]+tmp[65]*tmp[174]+tmp[66]*tmp[173]+tmp[67]*tmp[172]+tmp[68]*tmp[171]+tmp[69]*tmp[170]+tmp[70]*tmp[169]+tmp[71]*tmp[168]+tmp[72]*tmp[167]+tmp[73]*tmp[166]+tmp[74]*tmp[165]+tmp[75]*tmp[164]+tmp[76]*tmp[163]+tmp[77]*tmp[162]+tmp[78]*tmp[161]+tmp[79]*tmp[160]+tmp[80]*tmp[159]+tmp[81]*tmp[158]+tmp[82]*tmp[157]+tmp[83]*tmp[156]+tmp[84]*tmp[155]+tmp[85]*tmp[154]+tmp[86]*tmp[153]+tmp[87]*tmp[152]+tmp[88]*tmp[151]+tmp[89]*tmp[150]+tmp[90]*tmp[149]+tmp[91]*tmp[148]+tmp[92]*tmp[147]+tmp[93]*tmp[146]+tmp[94]*tmp[145]+tmp[95]*tmp[144]+tmp[96]*tmp[143]+tmp[97]*tmp[142]+tmp[98]*tmp[141]+tmp[99]*tmp[140];
				ans[140]<=tmp[41]*tmp[199]+tmp[42]*tmp[198]+tmp[43]*tmp[197]+tmp[44]*tmp[196]+tmp[45]*tmp[195]+tmp[46]*tmp[194]+tmp[47]*tmp[193]+tmp[48]*tmp[192]+tmp[49]*tmp[191]+tmp[50]*tmp[190]+tmp[51]*tmp[189]+tmp[52]*tmp[188]+tmp[53]*tmp[187]+tmp[54]*tmp[186]+tmp[55]*tmp[185]+tmp[56]*tmp[184]+tmp[57]*tmp[183]+tmp[58]*tmp[182]+tmp[59]*tmp[181]+tmp[60]*tmp[180]+tmp[61]*tmp[179]+tmp[62]*tmp[178]+tmp[63]*tmp[177]+tmp[64]*tmp[176]+tmp[65]*tmp[175]+tmp[66]*tmp[174]+tmp[67]*tmp[173]+tmp[68]*tmp[172]+tmp[69]*tmp[171]+tmp[70]*tmp[170]+tmp[71]*tmp[169]+tmp[72]*tmp[168]+tmp[73]*tmp[167]+tmp[74]*tmp[166]+tmp[75]*tmp[165]+tmp[76]*tmp[164]+tmp[77]*tmp[163]+tmp[78]*tmp[162]+tmp[79]*tmp[161]+tmp[80]*tmp[160]+tmp[81]*tmp[159]+tmp[82]*tmp[158]+tmp[83]*tmp[157]+tmp[84]*tmp[156]+tmp[85]*tmp[155]+tmp[86]*tmp[154]+tmp[87]*tmp[153]+tmp[88]*tmp[152]+tmp[89]*tmp[151]+tmp[90]*tmp[150]+tmp[91]*tmp[149]+tmp[92]*tmp[148]+tmp[93]*tmp[147]+tmp[94]*tmp[146]+tmp[95]*tmp[145]+tmp[96]*tmp[144]+tmp[97]*tmp[143]+tmp[98]*tmp[142]+tmp[99]*tmp[141];
				ans[141]<=tmp[42]*tmp[199]+tmp[43]*tmp[198]+tmp[44]*tmp[197]+tmp[45]*tmp[196]+tmp[46]*tmp[195]+tmp[47]*tmp[194]+tmp[48]*tmp[193]+tmp[49]*tmp[192]+tmp[50]*tmp[191]+tmp[51]*tmp[190]+tmp[52]*tmp[189]+tmp[53]*tmp[188]+tmp[54]*tmp[187]+tmp[55]*tmp[186]+tmp[56]*tmp[185]+tmp[57]*tmp[184]+tmp[58]*tmp[183]+tmp[59]*tmp[182]+tmp[60]*tmp[181]+tmp[61]*tmp[180]+tmp[62]*tmp[179]+tmp[63]*tmp[178]+tmp[64]*tmp[177]+tmp[65]*tmp[176]+tmp[66]*tmp[175]+tmp[67]*tmp[174]+tmp[68]*tmp[173]+tmp[69]*tmp[172]+tmp[70]*tmp[171]+tmp[71]*tmp[170]+tmp[72]*tmp[169]+tmp[73]*tmp[168]+tmp[74]*tmp[167]+tmp[75]*tmp[166]+tmp[76]*tmp[165]+tmp[77]*tmp[164]+tmp[78]*tmp[163]+tmp[79]*tmp[162]+tmp[80]*tmp[161]+tmp[81]*tmp[160]+tmp[82]*tmp[159]+tmp[83]*tmp[158]+tmp[84]*tmp[157]+tmp[85]*tmp[156]+tmp[86]*tmp[155]+tmp[87]*tmp[154]+tmp[88]*tmp[153]+tmp[89]*tmp[152]+tmp[90]*tmp[151]+tmp[91]*tmp[150]+tmp[92]*tmp[149]+tmp[93]*tmp[148]+tmp[94]*tmp[147]+tmp[95]*tmp[146]+tmp[96]*tmp[145]+tmp[97]*tmp[144]+tmp[98]*tmp[143]+tmp[99]*tmp[142];
				ans[142]<=tmp[43]*tmp[199]+tmp[44]*tmp[198]+tmp[45]*tmp[197]+tmp[46]*tmp[196]+tmp[47]*tmp[195]+tmp[48]*tmp[194]+tmp[49]*tmp[193]+tmp[50]*tmp[192]+tmp[51]*tmp[191]+tmp[52]*tmp[190]+tmp[53]*tmp[189]+tmp[54]*tmp[188]+tmp[55]*tmp[187]+tmp[56]*tmp[186]+tmp[57]*tmp[185]+tmp[58]*tmp[184]+tmp[59]*tmp[183]+tmp[60]*tmp[182]+tmp[61]*tmp[181]+tmp[62]*tmp[180]+tmp[63]*tmp[179]+tmp[64]*tmp[178]+tmp[65]*tmp[177]+tmp[66]*tmp[176]+tmp[67]*tmp[175]+tmp[68]*tmp[174]+tmp[69]*tmp[173]+tmp[70]*tmp[172]+tmp[71]*tmp[171]+tmp[72]*tmp[170]+tmp[73]*tmp[169]+tmp[74]*tmp[168]+tmp[75]*tmp[167]+tmp[76]*tmp[166]+tmp[77]*tmp[165]+tmp[78]*tmp[164]+tmp[79]*tmp[163]+tmp[80]*tmp[162]+tmp[81]*tmp[161]+tmp[82]*tmp[160]+tmp[83]*tmp[159]+tmp[84]*tmp[158]+tmp[85]*tmp[157]+tmp[86]*tmp[156]+tmp[87]*tmp[155]+tmp[88]*tmp[154]+tmp[89]*tmp[153]+tmp[90]*tmp[152]+tmp[91]*tmp[151]+tmp[92]*tmp[150]+tmp[93]*tmp[149]+tmp[94]*tmp[148]+tmp[95]*tmp[147]+tmp[96]*tmp[146]+tmp[97]*tmp[145]+tmp[98]*tmp[144]+tmp[99]*tmp[143];
				ans[143]<=tmp[44]*tmp[199]+tmp[45]*tmp[198]+tmp[46]*tmp[197]+tmp[47]*tmp[196]+tmp[48]*tmp[195]+tmp[49]*tmp[194]+tmp[50]*tmp[193]+tmp[51]*tmp[192]+tmp[52]*tmp[191]+tmp[53]*tmp[190]+tmp[54]*tmp[189]+tmp[55]*tmp[188]+tmp[56]*tmp[187]+tmp[57]*tmp[186]+tmp[58]*tmp[185]+tmp[59]*tmp[184]+tmp[60]*tmp[183]+tmp[61]*tmp[182]+tmp[62]*tmp[181]+tmp[63]*tmp[180]+tmp[64]*tmp[179]+tmp[65]*tmp[178]+tmp[66]*tmp[177]+tmp[67]*tmp[176]+tmp[68]*tmp[175]+tmp[69]*tmp[174]+tmp[70]*tmp[173]+tmp[71]*tmp[172]+tmp[72]*tmp[171]+tmp[73]*tmp[170]+tmp[74]*tmp[169]+tmp[75]*tmp[168]+tmp[76]*tmp[167]+tmp[77]*tmp[166]+tmp[78]*tmp[165]+tmp[79]*tmp[164]+tmp[80]*tmp[163]+tmp[81]*tmp[162]+tmp[82]*tmp[161]+tmp[83]*tmp[160]+tmp[84]*tmp[159]+tmp[85]*tmp[158]+tmp[86]*tmp[157]+tmp[87]*tmp[156]+tmp[88]*tmp[155]+tmp[89]*tmp[154]+tmp[90]*tmp[153]+tmp[91]*tmp[152]+tmp[92]*tmp[151]+tmp[93]*tmp[150]+tmp[94]*tmp[149]+tmp[95]*tmp[148]+tmp[96]*tmp[147]+tmp[97]*tmp[146]+tmp[98]*tmp[145]+tmp[99]*tmp[144];
				ans[144]<=tmp[45]*tmp[199]+tmp[46]*tmp[198]+tmp[47]*tmp[197]+tmp[48]*tmp[196]+tmp[49]*tmp[195]+tmp[50]*tmp[194]+tmp[51]*tmp[193]+tmp[52]*tmp[192]+tmp[53]*tmp[191]+tmp[54]*tmp[190]+tmp[55]*tmp[189]+tmp[56]*tmp[188]+tmp[57]*tmp[187]+tmp[58]*tmp[186]+tmp[59]*tmp[185]+tmp[60]*tmp[184]+tmp[61]*tmp[183]+tmp[62]*tmp[182]+tmp[63]*tmp[181]+tmp[64]*tmp[180]+tmp[65]*tmp[179]+tmp[66]*tmp[178]+tmp[67]*tmp[177]+tmp[68]*tmp[176]+tmp[69]*tmp[175]+tmp[70]*tmp[174]+tmp[71]*tmp[173]+tmp[72]*tmp[172]+tmp[73]*tmp[171]+tmp[74]*tmp[170]+tmp[75]*tmp[169]+tmp[76]*tmp[168]+tmp[77]*tmp[167]+tmp[78]*tmp[166]+tmp[79]*tmp[165]+tmp[80]*tmp[164]+tmp[81]*tmp[163]+tmp[82]*tmp[162]+tmp[83]*tmp[161]+tmp[84]*tmp[160]+tmp[85]*tmp[159]+tmp[86]*tmp[158]+tmp[87]*tmp[157]+tmp[88]*tmp[156]+tmp[89]*tmp[155]+tmp[90]*tmp[154]+tmp[91]*tmp[153]+tmp[92]*tmp[152]+tmp[93]*tmp[151]+tmp[94]*tmp[150]+tmp[95]*tmp[149]+tmp[96]*tmp[148]+tmp[97]*tmp[147]+tmp[98]*tmp[146]+tmp[99]*tmp[145];
				ans[145]<=tmp[46]*tmp[199]+tmp[47]*tmp[198]+tmp[48]*tmp[197]+tmp[49]*tmp[196]+tmp[50]*tmp[195]+tmp[51]*tmp[194]+tmp[52]*tmp[193]+tmp[53]*tmp[192]+tmp[54]*tmp[191]+tmp[55]*tmp[190]+tmp[56]*tmp[189]+tmp[57]*tmp[188]+tmp[58]*tmp[187]+tmp[59]*tmp[186]+tmp[60]*tmp[185]+tmp[61]*tmp[184]+tmp[62]*tmp[183]+tmp[63]*tmp[182]+tmp[64]*tmp[181]+tmp[65]*tmp[180]+tmp[66]*tmp[179]+tmp[67]*tmp[178]+tmp[68]*tmp[177]+tmp[69]*tmp[176]+tmp[70]*tmp[175]+tmp[71]*tmp[174]+tmp[72]*tmp[173]+tmp[73]*tmp[172]+tmp[74]*tmp[171]+tmp[75]*tmp[170]+tmp[76]*tmp[169]+tmp[77]*tmp[168]+tmp[78]*tmp[167]+tmp[79]*tmp[166]+tmp[80]*tmp[165]+tmp[81]*tmp[164]+tmp[82]*tmp[163]+tmp[83]*tmp[162]+tmp[84]*tmp[161]+tmp[85]*tmp[160]+tmp[86]*tmp[159]+tmp[87]*tmp[158]+tmp[88]*tmp[157]+tmp[89]*tmp[156]+tmp[90]*tmp[155]+tmp[91]*tmp[154]+tmp[92]*tmp[153]+tmp[93]*tmp[152]+tmp[94]*tmp[151]+tmp[95]*tmp[150]+tmp[96]*tmp[149]+tmp[97]*tmp[148]+tmp[98]*tmp[147]+tmp[99]*tmp[146];
				ans[146]<=tmp[47]*tmp[199]+tmp[48]*tmp[198]+tmp[49]*tmp[197]+tmp[50]*tmp[196]+tmp[51]*tmp[195]+tmp[52]*tmp[194]+tmp[53]*tmp[193]+tmp[54]*tmp[192]+tmp[55]*tmp[191]+tmp[56]*tmp[190]+tmp[57]*tmp[189]+tmp[58]*tmp[188]+tmp[59]*tmp[187]+tmp[60]*tmp[186]+tmp[61]*tmp[185]+tmp[62]*tmp[184]+tmp[63]*tmp[183]+tmp[64]*tmp[182]+tmp[65]*tmp[181]+tmp[66]*tmp[180]+tmp[67]*tmp[179]+tmp[68]*tmp[178]+tmp[69]*tmp[177]+tmp[70]*tmp[176]+tmp[71]*tmp[175]+tmp[72]*tmp[174]+tmp[73]*tmp[173]+tmp[74]*tmp[172]+tmp[75]*tmp[171]+tmp[76]*tmp[170]+tmp[77]*tmp[169]+tmp[78]*tmp[168]+tmp[79]*tmp[167]+tmp[80]*tmp[166]+tmp[81]*tmp[165]+tmp[82]*tmp[164]+tmp[83]*tmp[163]+tmp[84]*tmp[162]+tmp[85]*tmp[161]+tmp[86]*tmp[160]+tmp[87]*tmp[159]+tmp[88]*tmp[158]+tmp[89]*tmp[157]+tmp[90]*tmp[156]+tmp[91]*tmp[155]+tmp[92]*tmp[154]+tmp[93]*tmp[153]+tmp[94]*tmp[152]+tmp[95]*tmp[151]+tmp[96]*tmp[150]+tmp[97]*tmp[149]+tmp[98]*tmp[148]+tmp[99]*tmp[147];
				ans[147]<=tmp[48]*tmp[199]+tmp[49]*tmp[198]+tmp[50]*tmp[197]+tmp[51]*tmp[196]+tmp[52]*tmp[195]+tmp[53]*tmp[194]+tmp[54]*tmp[193]+tmp[55]*tmp[192]+tmp[56]*tmp[191]+tmp[57]*tmp[190]+tmp[58]*tmp[189]+tmp[59]*tmp[188]+tmp[60]*tmp[187]+tmp[61]*tmp[186]+tmp[62]*tmp[185]+tmp[63]*tmp[184]+tmp[64]*tmp[183]+tmp[65]*tmp[182]+tmp[66]*tmp[181]+tmp[67]*tmp[180]+tmp[68]*tmp[179]+tmp[69]*tmp[178]+tmp[70]*tmp[177]+tmp[71]*tmp[176]+tmp[72]*tmp[175]+tmp[73]*tmp[174]+tmp[74]*tmp[173]+tmp[75]*tmp[172]+tmp[76]*tmp[171]+tmp[77]*tmp[170]+tmp[78]*tmp[169]+tmp[79]*tmp[168]+tmp[80]*tmp[167]+tmp[81]*tmp[166]+tmp[82]*tmp[165]+tmp[83]*tmp[164]+tmp[84]*tmp[163]+tmp[85]*tmp[162]+tmp[86]*tmp[161]+tmp[87]*tmp[160]+tmp[88]*tmp[159]+tmp[89]*tmp[158]+tmp[90]*tmp[157]+tmp[91]*tmp[156]+tmp[92]*tmp[155]+tmp[93]*tmp[154]+tmp[94]*tmp[153]+tmp[95]*tmp[152]+tmp[96]*tmp[151]+tmp[97]*tmp[150]+tmp[98]*tmp[149]+tmp[99]*tmp[148];
				ans[148]<=tmp[49]*tmp[199]+tmp[50]*tmp[198]+tmp[51]*tmp[197]+tmp[52]*tmp[196]+tmp[53]*tmp[195]+tmp[54]*tmp[194]+tmp[55]*tmp[193]+tmp[56]*tmp[192]+tmp[57]*tmp[191]+tmp[58]*tmp[190]+tmp[59]*tmp[189]+tmp[60]*tmp[188]+tmp[61]*tmp[187]+tmp[62]*tmp[186]+tmp[63]*tmp[185]+tmp[64]*tmp[184]+tmp[65]*tmp[183]+tmp[66]*tmp[182]+tmp[67]*tmp[181]+tmp[68]*tmp[180]+tmp[69]*tmp[179]+tmp[70]*tmp[178]+tmp[71]*tmp[177]+tmp[72]*tmp[176]+tmp[73]*tmp[175]+tmp[74]*tmp[174]+tmp[75]*tmp[173]+tmp[76]*tmp[172]+tmp[77]*tmp[171]+tmp[78]*tmp[170]+tmp[79]*tmp[169]+tmp[80]*tmp[168]+tmp[81]*tmp[167]+tmp[82]*tmp[166]+tmp[83]*tmp[165]+tmp[84]*tmp[164]+tmp[85]*tmp[163]+tmp[86]*tmp[162]+tmp[87]*tmp[161]+tmp[88]*tmp[160]+tmp[89]*tmp[159]+tmp[90]*tmp[158]+tmp[91]*tmp[157]+tmp[92]*tmp[156]+tmp[93]*tmp[155]+tmp[94]*tmp[154]+tmp[95]*tmp[153]+tmp[96]*tmp[152]+tmp[97]*tmp[151]+tmp[98]*tmp[150]+tmp[99]*tmp[149];
				ans[149]<=tmp[50]*tmp[199]+tmp[51]*tmp[198]+tmp[52]*tmp[197]+tmp[53]*tmp[196]+tmp[54]*tmp[195]+tmp[55]*tmp[194]+tmp[56]*tmp[193]+tmp[57]*tmp[192]+tmp[58]*tmp[191]+tmp[59]*tmp[190]+tmp[60]*tmp[189]+tmp[61]*tmp[188]+tmp[62]*tmp[187]+tmp[63]*tmp[186]+tmp[64]*tmp[185]+tmp[65]*tmp[184]+tmp[66]*tmp[183]+tmp[67]*tmp[182]+tmp[68]*tmp[181]+tmp[69]*tmp[180]+tmp[70]*tmp[179]+tmp[71]*tmp[178]+tmp[72]*tmp[177]+tmp[73]*tmp[176]+tmp[74]*tmp[175]+tmp[75]*tmp[174]+tmp[76]*tmp[173]+tmp[77]*tmp[172]+tmp[78]*tmp[171]+tmp[79]*tmp[170]+tmp[80]*tmp[169]+tmp[81]*tmp[168]+tmp[82]*tmp[167]+tmp[83]*tmp[166]+tmp[84]*tmp[165]+tmp[85]*tmp[164]+tmp[86]*tmp[163]+tmp[87]*tmp[162]+tmp[88]*tmp[161]+tmp[89]*tmp[160]+tmp[90]*tmp[159]+tmp[91]*tmp[158]+tmp[92]*tmp[157]+tmp[93]*tmp[156]+tmp[94]*tmp[155]+tmp[95]*tmp[154]+tmp[96]*tmp[153]+tmp[97]*tmp[152]+tmp[98]*tmp[151]+tmp[99]*tmp[150];
				ans[150]<=tmp[51]*tmp[199]+tmp[52]*tmp[198]+tmp[53]*tmp[197]+tmp[54]*tmp[196]+tmp[55]*tmp[195]+tmp[56]*tmp[194]+tmp[57]*tmp[193]+tmp[58]*tmp[192]+tmp[59]*tmp[191]+tmp[60]*tmp[190]+tmp[61]*tmp[189]+tmp[62]*tmp[188]+tmp[63]*tmp[187]+tmp[64]*tmp[186]+tmp[65]*tmp[185]+tmp[66]*tmp[184]+tmp[67]*tmp[183]+tmp[68]*tmp[182]+tmp[69]*tmp[181]+tmp[70]*tmp[180]+tmp[71]*tmp[179]+tmp[72]*tmp[178]+tmp[73]*tmp[177]+tmp[74]*tmp[176]+tmp[75]*tmp[175]+tmp[76]*tmp[174]+tmp[77]*tmp[173]+tmp[78]*tmp[172]+tmp[79]*tmp[171]+tmp[80]*tmp[170]+tmp[81]*tmp[169]+tmp[82]*tmp[168]+tmp[83]*tmp[167]+tmp[84]*tmp[166]+tmp[85]*tmp[165]+tmp[86]*tmp[164]+tmp[87]*tmp[163]+tmp[88]*tmp[162]+tmp[89]*tmp[161]+tmp[90]*tmp[160]+tmp[91]*tmp[159]+tmp[92]*tmp[158]+tmp[93]*tmp[157]+tmp[94]*tmp[156]+tmp[95]*tmp[155]+tmp[96]*tmp[154]+tmp[97]*tmp[153]+tmp[98]*tmp[152]+tmp[99]*tmp[151];
				ans[151]<=tmp[52]*tmp[199]+tmp[53]*tmp[198]+tmp[54]*tmp[197]+tmp[55]*tmp[196]+tmp[56]*tmp[195]+tmp[57]*tmp[194]+tmp[58]*tmp[193]+tmp[59]*tmp[192]+tmp[60]*tmp[191]+tmp[61]*tmp[190]+tmp[62]*tmp[189]+tmp[63]*tmp[188]+tmp[64]*tmp[187]+tmp[65]*tmp[186]+tmp[66]*tmp[185]+tmp[67]*tmp[184]+tmp[68]*tmp[183]+tmp[69]*tmp[182]+tmp[70]*tmp[181]+tmp[71]*tmp[180]+tmp[72]*tmp[179]+tmp[73]*tmp[178]+tmp[74]*tmp[177]+tmp[75]*tmp[176]+tmp[76]*tmp[175]+tmp[77]*tmp[174]+tmp[78]*tmp[173]+tmp[79]*tmp[172]+tmp[80]*tmp[171]+tmp[81]*tmp[170]+tmp[82]*tmp[169]+tmp[83]*tmp[168]+tmp[84]*tmp[167]+tmp[85]*tmp[166]+tmp[86]*tmp[165]+tmp[87]*tmp[164]+tmp[88]*tmp[163]+tmp[89]*tmp[162]+tmp[90]*tmp[161]+tmp[91]*tmp[160]+tmp[92]*tmp[159]+tmp[93]*tmp[158]+tmp[94]*tmp[157]+tmp[95]*tmp[156]+tmp[96]*tmp[155]+tmp[97]*tmp[154]+tmp[98]*tmp[153]+tmp[99]*tmp[152];
				ans[152]<=tmp[53]*tmp[199]+tmp[54]*tmp[198]+tmp[55]*tmp[197]+tmp[56]*tmp[196]+tmp[57]*tmp[195]+tmp[58]*tmp[194]+tmp[59]*tmp[193]+tmp[60]*tmp[192]+tmp[61]*tmp[191]+tmp[62]*tmp[190]+tmp[63]*tmp[189]+tmp[64]*tmp[188]+tmp[65]*tmp[187]+tmp[66]*tmp[186]+tmp[67]*tmp[185]+tmp[68]*tmp[184]+tmp[69]*tmp[183]+tmp[70]*tmp[182]+tmp[71]*tmp[181]+tmp[72]*tmp[180]+tmp[73]*tmp[179]+tmp[74]*tmp[178]+tmp[75]*tmp[177]+tmp[76]*tmp[176]+tmp[77]*tmp[175]+tmp[78]*tmp[174]+tmp[79]*tmp[173]+tmp[80]*tmp[172]+tmp[81]*tmp[171]+tmp[82]*tmp[170]+tmp[83]*tmp[169]+tmp[84]*tmp[168]+tmp[85]*tmp[167]+tmp[86]*tmp[166]+tmp[87]*tmp[165]+tmp[88]*tmp[164]+tmp[89]*tmp[163]+tmp[90]*tmp[162]+tmp[91]*tmp[161]+tmp[92]*tmp[160]+tmp[93]*tmp[159]+tmp[94]*tmp[158]+tmp[95]*tmp[157]+tmp[96]*tmp[156]+tmp[97]*tmp[155]+tmp[98]*tmp[154]+tmp[99]*tmp[153];
				ans[153]<=tmp[54]*tmp[199]+tmp[55]*tmp[198]+tmp[56]*tmp[197]+tmp[57]*tmp[196]+tmp[58]*tmp[195]+tmp[59]*tmp[194]+tmp[60]*tmp[193]+tmp[61]*tmp[192]+tmp[62]*tmp[191]+tmp[63]*tmp[190]+tmp[64]*tmp[189]+tmp[65]*tmp[188]+tmp[66]*tmp[187]+tmp[67]*tmp[186]+tmp[68]*tmp[185]+tmp[69]*tmp[184]+tmp[70]*tmp[183]+tmp[71]*tmp[182]+tmp[72]*tmp[181]+tmp[73]*tmp[180]+tmp[74]*tmp[179]+tmp[75]*tmp[178]+tmp[76]*tmp[177]+tmp[77]*tmp[176]+tmp[78]*tmp[175]+tmp[79]*tmp[174]+tmp[80]*tmp[173]+tmp[81]*tmp[172]+tmp[82]*tmp[171]+tmp[83]*tmp[170]+tmp[84]*tmp[169]+tmp[85]*tmp[168]+tmp[86]*tmp[167]+tmp[87]*tmp[166]+tmp[88]*tmp[165]+tmp[89]*tmp[164]+tmp[90]*tmp[163]+tmp[91]*tmp[162]+tmp[92]*tmp[161]+tmp[93]*tmp[160]+tmp[94]*tmp[159]+tmp[95]*tmp[158]+tmp[96]*tmp[157]+tmp[97]*tmp[156]+tmp[98]*tmp[155]+tmp[99]*tmp[154];
				ans[154]<=tmp[55]*tmp[199]+tmp[56]*tmp[198]+tmp[57]*tmp[197]+tmp[58]*tmp[196]+tmp[59]*tmp[195]+tmp[60]*tmp[194]+tmp[61]*tmp[193]+tmp[62]*tmp[192]+tmp[63]*tmp[191]+tmp[64]*tmp[190]+tmp[65]*tmp[189]+tmp[66]*tmp[188]+tmp[67]*tmp[187]+tmp[68]*tmp[186]+tmp[69]*tmp[185]+tmp[70]*tmp[184]+tmp[71]*tmp[183]+tmp[72]*tmp[182]+tmp[73]*tmp[181]+tmp[74]*tmp[180]+tmp[75]*tmp[179]+tmp[76]*tmp[178]+tmp[77]*tmp[177]+tmp[78]*tmp[176]+tmp[79]*tmp[175]+tmp[80]*tmp[174]+tmp[81]*tmp[173]+tmp[82]*tmp[172]+tmp[83]*tmp[171]+tmp[84]*tmp[170]+tmp[85]*tmp[169]+tmp[86]*tmp[168]+tmp[87]*tmp[167]+tmp[88]*tmp[166]+tmp[89]*tmp[165]+tmp[90]*tmp[164]+tmp[91]*tmp[163]+tmp[92]*tmp[162]+tmp[93]*tmp[161]+tmp[94]*tmp[160]+tmp[95]*tmp[159]+tmp[96]*tmp[158]+tmp[97]*tmp[157]+tmp[98]*tmp[156]+tmp[99]*tmp[155];
				ans[155]<=tmp[56]*tmp[199]+tmp[57]*tmp[198]+tmp[58]*tmp[197]+tmp[59]*tmp[196]+tmp[60]*tmp[195]+tmp[61]*tmp[194]+tmp[62]*tmp[193]+tmp[63]*tmp[192]+tmp[64]*tmp[191]+tmp[65]*tmp[190]+tmp[66]*tmp[189]+tmp[67]*tmp[188]+tmp[68]*tmp[187]+tmp[69]*tmp[186]+tmp[70]*tmp[185]+tmp[71]*tmp[184]+tmp[72]*tmp[183]+tmp[73]*tmp[182]+tmp[74]*tmp[181]+tmp[75]*tmp[180]+tmp[76]*tmp[179]+tmp[77]*tmp[178]+tmp[78]*tmp[177]+tmp[79]*tmp[176]+tmp[80]*tmp[175]+tmp[81]*tmp[174]+tmp[82]*tmp[173]+tmp[83]*tmp[172]+tmp[84]*tmp[171]+tmp[85]*tmp[170]+tmp[86]*tmp[169]+tmp[87]*tmp[168]+tmp[88]*tmp[167]+tmp[89]*tmp[166]+tmp[90]*tmp[165]+tmp[91]*tmp[164]+tmp[92]*tmp[163]+tmp[93]*tmp[162]+tmp[94]*tmp[161]+tmp[95]*tmp[160]+tmp[96]*tmp[159]+tmp[97]*tmp[158]+tmp[98]*tmp[157]+tmp[99]*tmp[156];
				ans[156]<=tmp[57]*tmp[199]+tmp[58]*tmp[198]+tmp[59]*tmp[197]+tmp[60]*tmp[196]+tmp[61]*tmp[195]+tmp[62]*tmp[194]+tmp[63]*tmp[193]+tmp[64]*tmp[192]+tmp[65]*tmp[191]+tmp[66]*tmp[190]+tmp[67]*tmp[189]+tmp[68]*tmp[188]+tmp[69]*tmp[187]+tmp[70]*tmp[186]+tmp[71]*tmp[185]+tmp[72]*tmp[184]+tmp[73]*tmp[183]+tmp[74]*tmp[182]+tmp[75]*tmp[181]+tmp[76]*tmp[180]+tmp[77]*tmp[179]+tmp[78]*tmp[178]+tmp[79]*tmp[177]+tmp[80]*tmp[176]+tmp[81]*tmp[175]+tmp[82]*tmp[174]+tmp[83]*tmp[173]+tmp[84]*tmp[172]+tmp[85]*tmp[171]+tmp[86]*tmp[170]+tmp[87]*tmp[169]+tmp[88]*tmp[168]+tmp[89]*tmp[167]+tmp[90]*tmp[166]+tmp[91]*tmp[165]+tmp[92]*tmp[164]+tmp[93]*tmp[163]+tmp[94]*tmp[162]+tmp[95]*tmp[161]+tmp[96]*tmp[160]+tmp[97]*tmp[159]+tmp[98]*tmp[158]+tmp[99]*tmp[157];
				ans[157]<=tmp[58]*tmp[199]+tmp[59]*tmp[198]+tmp[60]*tmp[197]+tmp[61]*tmp[196]+tmp[62]*tmp[195]+tmp[63]*tmp[194]+tmp[64]*tmp[193]+tmp[65]*tmp[192]+tmp[66]*tmp[191]+tmp[67]*tmp[190]+tmp[68]*tmp[189]+tmp[69]*tmp[188]+tmp[70]*tmp[187]+tmp[71]*tmp[186]+tmp[72]*tmp[185]+tmp[73]*tmp[184]+tmp[74]*tmp[183]+tmp[75]*tmp[182]+tmp[76]*tmp[181]+tmp[77]*tmp[180]+tmp[78]*tmp[179]+tmp[79]*tmp[178]+tmp[80]*tmp[177]+tmp[81]*tmp[176]+tmp[82]*tmp[175]+tmp[83]*tmp[174]+tmp[84]*tmp[173]+tmp[85]*tmp[172]+tmp[86]*tmp[171]+tmp[87]*tmp[170]+tmp[88]*tmp[169]+tmp[89]*tmp[168]+tmp[90]*tmp[167]+tmp[91]*tmp[166]+tmp[92]*tmp[165]+tmp[93]*tmp[164]+tmp[94]*tmp[163]+tmp[95]*tmp[162]+tmp[96]*tmp[161]+tmp[97]*tmp[160]+tmp[98]*tmp[159]+tmp[99]*tmp[158];
				ans[158]<=tmp[59]*tmp[199]+tmp[60]*tmp[198]+tmp[61]*tmp[197]+tmp[62]*tmp[196]+tmp[63]*tmp[195]+tmp[64]*tmp[194]+tmp[65]*tmp[193]+tmp[66]*tmp[192]+tmp[67]*tmp[191]+tmp[68]*tmp[190]+tmp[69]*tmp[189]+tmp[70]*tmp[188]+tmp[71]*tmp[187]+tmp[72]*tmp[186]+tmp[73]*tmp[185]+tmp[74]*tmp[184]+tmp[75]*tmp[183]+tmp[76]*tmp[182]+tmp[77]*tmp[181]+tmp[78]*tmp[180]+tmp[79]*tmp[179]+tmp[80]*tmp[178]+tmp[81]*tmp[177]+tmp[82]*tmp[176]+tmp[83]*tmp[175]+tmp[84]*tmp[174]+tmp[85]*tmp[173]+tmp[86]*tmp[172]+tmp[87]*tmp[171]+tmp[88]*tmp[170]+tmp[89]*tmp[169]+tmp[90]*tmp[168]+tmp[91]*tmp[167]+tmp[92]*tmp[166]+tmp[93]*tmp[165]+tmp[94]*tmp[164]+tmp[95]*tmp[163]+tmp[96]*tmp[162]+tmp[97]*tmp[161]+tmp[98]*tmp[160]+tmp[99]*tmp[159];
				ans[159]<=tmp[60]*tmp[199]+tmp[61]*tmp[198]+tmp[62]*tmp[197]+tmp[63]*tmp[196]+tmp[64]*tmp[195]+tmp[65]*tmp[194]+tmp[66]*tmp[193]+tmp[67]*tmp[192]+tmp[68]*tmp[191]+tmp[69]*tmp[190]+tmp[70]*tmp[189]+tmp[71]*tmp[188]+tmp[72]*tmp[187]+tmp[73]*tmp[186]+tmp[74]*tmp[185]+tmp[75]*tmp[184]+tmp[76]*tmp[183]+tmp[77]*tmp[182]+tmp[78]*tmp[181]+tmp[79]*tmp[180]+tmp[80]*tmp[179]+tmp[81]*tmp[178]+tmp[82]*tmp[177]+tmp[83]*tmp[176]+tmp[84]*tmp[175]+tmp[85]*tmp[174]+tmp[86]*tmp[173]+tmp[87]*tmp[172]+tmp[88]*tmp[171]+tmp[89]*tmp[170]+tmp[90]*tmp[169]+tmp[91]*tmp[168]+tmp[92]*tmp[167]+tmp[93]*tmp[166]+tmp[94]*tmp[165]+tmp[95]*tmp[164]+tmp[96]*tmp[163]+tmp[97]*tmp[162]+tmp[98]*tmp[161]+tmp[99]*tmp[160];
				ans[160]<=tmp[61]*tmp[199]+tmp[62]*tmp[198]+tmp[63]*tmp[197]+tmp[64]*tmp[196]+tmp[65]*tmp[195]+tmp[66]*tmp[194]+tmp[67]*tmp[193]+tmp[68]*tmp[192]+tmp[69]*tmp[191]+tmp[70]*tmp[190]+tmp[71]*tmp[189]+tmp[72]*tmp[188]+tmp[73]*tmp[187]+tmp[74]*tmp[186]+tmp[75]*tmp[185]+tmp[76]*tmp[184]+tmp[77]*tmp[183]+tmp[78]*tmp[182]+tmp[79]*tmp[181]+tmp[80]*tmp[180]+tmp[81]*tmp[179]+tmp[82]*tmp[178]+tmp[83]*tmp[177]+tmp[84]*tmp[176]+tmp[85]*tmp[175]+tmp[86]*tmp[174]+tmp[87]*tmp[173]+tmp[88]*tmp[172]+tmp[89]*tmp[171]+tmp[90]*tmp[170]+tmp[91]*tmp[169]+tmp[92]*tmp[168]+tmp[93]*tmp[167]+tmp[94]*tmp[166]+tmp[95]*tmp[165]+tmp[96]*tmp[164]+tmp[97]*tmp[163]+tmp[98]*tmp[162]+tmp[99]*tmp[161];
				ans[161]<=tmp[62]*tmp[199]+tmp[63]*tmp[198]+tmp[64]*tmp[197]+tmp[65]*tmp[196]+tmp[66]*tmp[195]+tmp[67]*tmp[194]+tmp[68]*tmp[193]+tmp[69]*tmp[192]+tmp[70]*tmp[191]+tmp[71]*tmp[190]+tmp[72]*tmp[189]+tmp[73]*tmp[188]+tmp[74]*tmp[187]+tmp[75]*tmp[186]+tmp[76]*tmp[185]+tmp[77]*tmp[184]+tmp[78]*tmp[183]+tmp[79]*tmp[182]+tmp[80]*tmp[181]+tmp[81]*tmp[180]+tmp[82]*tmp[179]+tmp[83]*tmp[178]+tmp[84]*tmp[177]+tmp[85]*tmp[176]+tmp[86]*tmp[175]+tmp[87]*tmp[174]+tmp[88]*tmp[173]+tmp[89]*tmp[172]+tmp[90]*tmp[171]+tmp[91]*tmp[170]+tmp[92]*tmp[169]+tmp[93]*tmp[168]+tmp[94]*tmp[167]+tmp[95]*tmp[166]+tmp[96]*tmp[165]+tmp[97]*tmp[164]+tmp[98]*tmp[163]+tmp[99]*tmp[162];
				ans[162]<=tmp[63]*tmp[199]+tmp[64]*tmp[198]+tmp[65]*tmp[197]+tmp[66]*tmp[196]+tmp[67]*tmp[195]+tmp[68]*tmp[194]+tmp[69]*tmp[193]+tmp[70]*tmp[192]+tmp[71]*tmp[191]+tmp[72]*tmp[190]+tmp[73]*tmp[189]+tmp[74]*tmp[188]+tmp[75]*tmp[187]+tmp[76]*tmp[186]+tmp[77]*tmp[185]+tmp[78]*tmp[184]+tmp[79]*tmp[183]+tmp[80]*tmp[182]+tmp[81]*tmp[181]+tmp[82]*tmp[180]+tmp[83]*tmp[179]+tmp[84]*tmp[178]+tmp[85]*tmp[177]+tmp[86]*tmp[176]+tmp[87]*tmp[175]+tmp[88]*tmp[174]+tmp[89]*tmp[173]+tmp[90]*tmp[172]+tmp[91]*tmp[171]+tmp[92]*tmp[170]+tmp[93]*tmp[169]+tmp[94]*tmp[168]+tmp[95]*tmp[167]+tmp[96]*tmp[166]+tmp[97]*tmp[165]+tmp[98]*tmp[164]+tmp[99]*tmp[163];
				ans[163]<=tmp[64]*tmp[199]+tmp[65]*tmp[198]+tmp[66]*tmp[197]+tmp[67]*tmp[196]+tmp[68]*tmp[195]+tmp[69]*tmp[194]+tmp[70]*tmp[193]+tmp[71]*tmp[192]+tmp[72]*tmp[191]+tmp[73]*tmp[190]+tmp[74]*tmp[189]+tmp[75]*tmp[188]+tmp[76]*tmp[187]+tmp[77]*tmp[186]+tmp[78]*tmp[185]+tmp[79]*tmp[184]+tmp[80]*tmp[183]+tmp[81]*tmp[182]+tmp[82]*tmp[181]+tmp[83]*tmp[180]+tmp[84]*tmp[179]+tmp[85]*tmp[178]+tmp[86]*tmp[177]+tmp[87]*tmp[176]+tmp[88]*tmp[175]+tmp[89]*tmp[174]+tmp[90]*tmp[173]+tmp[91]*tmp[172]+tmp[92]*tmp[171]+tmp[93]*tmp[170]+tmp[94]*tmp[169]+tmp[95]*tmp[168]+tmp[96]*tmp[167]+tmp[97]*tmp[166]+tmp[98]*tmp[165]+tmp[99]*tmp[164];
				ans[164]<=tmp[65]*tmp[199]+tmp[66]*tmp[198]+tmp[67]*tmp[197]+tmp[68]*tmp[196]+tmp[69]*tmp[195]+tmp[70]*tmp[194]+tmp[71]*tmp[193]+tmp[72]*tmp[192]+tmp[73]*tmp[191]+tmp[74]*tmp[190]+tmp[75]*tmp[189]+tmp[76]*tmp[188]+tmp[77]*tmp[187]+tmp[78]*tmp[186]+tmp[79]*tmp[185]+tmp[80]*tmp[184]+tmp[81]*tmp[183]+tmp[82]*tmp[182]+tmp[83]*tmp[181]+tmp[84]*tmp[180]+tmp[85]*tmp[179]+tmp[86]*tmp[178]+tmp[87]*tmp[177]+tmp[88]*tmp[176]+tmp[89]*tmp[175]+tmp[90]*tmp[174]+tmp[91]*tmp[173]+tmp[92]*tmp[172]+tmp[93]*tmp[171]+tmp[94]*tmp[170]+tmp[95]*tmp[169]+tmp[96]*tmp[168]+tmp[97]*tmp[167]+tmp[98]*tmp[166]+tmp[99]*tmp[165];
				ans[165]<=tmp[66]*tmp[199]+tmp[67]*tmp[198]+tmp[68]*tmp[197]+tmp[69]*tmp[196]+tmp[70]*tmp[195]+tmp[71]*tmp[194]+tmp[72]*tmp[193]+tmp[73]*tmp[192]+tmp[74]*tmp[191]+tmp[75]*tmp[190]+tmp[76]*tmp[189]+tmp[77]*tmp[188]+tmp[78]*tmp[187]+tmp[79]*tmp[186]+tmp[80]*tmp[185]+tmp[81]*tmp[184]+tmp[82]*tmp[183]+tmp[83]*tmp[182]+tmp[84]*tmp[181]+tmp[85]*tmp[180]+tmp[86]*tmp[179]+tmp[87]*tmp[178]+tmp[88]*tmp[177]+tmp[89]*tmp[176]+tmp[90]*tmp[175]+tmp[91]*tmp[174]+tmp[92]*tmp[173]+tmp[93]*tmp[172]+tmp[94]*tmp[171]+tmp[95]*tmp[170]+tmp[96]*tmp[169]+tmp[97]*tmp[168]+tmp[98]*tmp[167]+tmp[99]*tmp[166];
				ans[166]<=tmp[67]*tmp[199]+tmp[68]*tmp[198]+tmp[69]*tmp[197]+tmp[70]*tmp[196]+tmp[71]*tmp[195]+tmp[72]*tmp[194]+tmp[73]*tmp[193]+tmp[74]*tmp[192]+tmp[75]*tmp[191]+tmp[76]*tmp[190]+tmp[77]*tmp[189]+tmp[78]*tmp[188]+tmp[79]*tmp[187]+tmp[80]*tmp[186]+tmp[81]*tmp[185]+tmp[82]*tmp[184]+tmp[83]*tmp[183]+tmp[84]*tmp[182]+tmp[85]*tmp[181]+tmp[86]*tmp[180]+tmp[87]*tmp[179]+tmp[88]*tmp[178]+tmp[89]*tmp[177]+tmp[90]*tmp[176]+tmp[91]*tmp[175]+tmp[92]*tmp[174]+tmp[93]*tmp[173]+tmp[94]*tmp[172]+tmp[95]*tmp[171]+tmp[96]*tmp[170]+tmp[97]*tmp[169]+tmp[98]*tmp[168]+tmp[99]*tmp[167];
				ans[167]<=tmp[68]*tmp[199]+tmp[69]*tmp[198]+tmp[70]*tmp[197]+tmp[71]*tmp[196]+tmp[72]*tmp[195]+tmp[73]*tmp[194]+tmp[74]*tmp[193]+tmp[75]*tmp[192]+tmp[76]*tmp[191]+tmp[77]*tmp[190]+tmp[78]*tmp[189]+tmp[79]*tmp[188]+tmp[80]*tmp[187]+tmp[81]*tmp[186]+tmp[82]*tmp[185]+tmp[83]*tmp[184]+tmp[84]*tmp[183]+tmp[85]*tmp[182]+tmp[86]*tmp[181]+tmp[87]*tmp[180]+tmp[88]*tmp[179]+tmp[89]*tmp[178]+tmp[90]*tmp[177]+tmp[91]*tmp[176]+tmp[92]*tmp[175]+tmp[93]*tmp[174]+tmp[94]*tmp[173]+tmp[95]*tmp[172]+tmp[96]*tmp[171]+tmp[97]*tmp[170]+tmp[98]*tmp[169]+tmp[99]*tmp[168];
				ans[168]<=tmp[69]*tmp[199]+tmp[70]*tmp[198]+tmp[71]*tmp[197]+tmp[72]*tmp[196]+tmp[73]*tmp[195]+tmp[74]*tmp[194]+tmp[75]*tmp[193]+tmp[76]*tmp[192]+tmp[77]*tmp[191]+tmp[78]*tmp[190]+tmp[79]*tmp[189]+tmp[80]*tmp[188]+tmp[81]*tmp[187]+tmp[82]*tmp[186]+tmp[83]*tmp[185]+tmp[84]*tmp[184]+tmp[85]*tmp[183]+tmp[86]*tmp[182]+tmp[87]*tmp[181]+tmp[88]*tmp[180]+tmp[89]*tmp[179]+tmp[90]*tmp[178]+tmp[91]*tmp[177]+tmp[92]*tmp[176]+tmp[93]*tmp[175]+tmp[94]*tmp[174]+tmp[95]*tmp[173]+tmp[96]*tmp[172]+tmp[97]*tmp[171]+tmp[98]*tmp[170]+tmp[99]*tmp[169];
				ans[169]<=tmp[70]*tmp[199]+tmp[71]*tmp[198]+tmp[72]*tmp[197]+tmp[73]*tmp[196]+tmp[74]*tmp[195]+tmp[75]*tmp[194]+tmp[76]*tmp[193]+tmp[77]*tmp[192]+tmp[78]*tmp[191]+tmp[79]*tmp[190]+tmp[80]*tmp[189]+tmp[81]*tmp[188]+tmp[82]*tmp[187]+tmp[83]*tmp[186]+tmp[84]*tmp[185]+tmp[85]*tmp[184]+tmp[86]*tmp[183]+tmp[87]*tmp[182]+tmp[88]*tmp[181]+tmp[89]*tmp[180]+tmp[90]*tmp[179]+tmp[91]*tmp[178]+tmp[92]*tmp[177]+tmp[93]*tmp[176]+tmp[94]*tmp[175]+tmp[95]*tmp[174]+tmp[96]*tmp[173]+tmp[97]*tmp[172]+tmp[98]*tmp[171]+tmp[99]*tmp[170];
				ans[170]<=tmp[71]*tmp[199]+tmp[72]*tmp[198]+tmp[73]*tmp[197]+tmp[74]*tmp[196]+tmp[75]*tmp[195]+tmp[76]*tmp[194]+tmp[77]*tmp[193]+tmp[78]*tmp[192]+tmp[79]*tmp[191]+tmp[80]*tmp[190]+tmp[81]*tmp[189]+tmp[82]*tmp[188]+tmp[83]*tmp[187]+tmp[84]*tmp[186]+tmp[85]*tmp[185]+tmp[86]*tmp[184]+tmp[87]*tmp[183]+tmp[88]*tmp[182]+tmp[89]*tmp[181]+tmp[90]*tmp[180]+tmp[91]*tmp[179]+tmp[92]*tmp[178]+tmp[93]*tmp[177]+tmp[94]*tmp[176]+tmp[95]*tmp[175]+tmp[96]*tmp[174]+tmp[97]*tmp[173]+tmp[98]*tmp[172]+tmp[99]*tmp[171];
				ans[171]<=tmp[72]*tmp[199]+tmp[73]*tmp[198]+tmp[74]*tmp[197]+tmp[75]*tmp[196]+tmp[76]*tmp[195]+tmp[77]*tmp[194]+tmp[78]*tmp[193]+tmp[79]*tmp[192]+tmp[80]*tmp[191]+tmp[81]*tmp[190]+tmp[82]*tmp[189]+tmp[83]*tmp[188]+tmp[84]*tmp[187]+tmp[85]*tmp[186]+tmp[86]*tmp[185]+tmp[87]*tmp[184]+tmp[88]*tmp[183]+tmp[89]*tmp[182]+tmp[90]*tmp[181]+tmp[91]*tmp[180]+tmp[92]*tmp[179]+tmp[93]*tmp[178]+tmp[94]*tmp[177]+tmp[95]*tmp[176]+tmp[96]*tmp[175]+tmp[97]*tmp[174]+tmp[98]*tmp[173]+tmp[99]*tmp[172];
				ans[172]<=tmp[73]*tmp[199]+tmp[74]*tmp[198]+tmp[75]*tmp[197]+tmp[76]*tmp[196]+tmp[77]*tmp[195]+tmp[78]*tmp[194]+tmp[79]*tmp[193]+tmp[80]*tmp[192]+tmp[81]*tmp[191]+tmp[82]*tmp[190]+tmp[83]*tmp[189]+tmp[84]*tmp[188]+tmp[85]*tmp[187]+tmp[86]*tmp[186]+tmp[87]*tmp[185]+tmp[88]*tmp[184]+tmp[89]*tmp[183]+tmp[90]*tmp[182]+tmp[91]*tmp[181]+tmp[92]*tmp[180]+tmp[93]*tmp[179]+tmp[94]*tmp[178]+tmp[95]*tmp[177]+tmp[96]*tmp[176]+tmp[97]*tmp[175]+tmp[98]*tmp[174]+tmp[99]*tmp[173];
				ans[173]<=tmp[74]*tmp[199]+tmp[75]*tmp[198]+tmp[76]*tmp[197]+tmp[77]*tmp[196]+tmp[78]*tmp[195]+tmp[79]*tmp[194]+tmp[80]*tmp[193]+tmp[81]*tmp[192]+tmp[82]*tmp[191]+tmp[83]*tmp[190]+tmp[84]*tmp[189]+tmp[85]*tmp[188]+tmp[86]*tmp[187]+tmp[87]*tmp[186]+tmp[88]*tmp[185]+tmp[89]*tmp[184]+tmp[90]*tmp[183]+tmp[91]*tmp[182]+tmp[92]*tmp[181]+tmp[93]*tmp[180]+tmp[94]*tmp[179]+tmp[95]*tmp[178]+tmp[96]*tmp[177]+tmp[97]*tmp[176]+tmp[98]*tmp[175]+tmp[99]*tmp[174];
				ans[174]<=tmp[75]*tmp[199]+tmp[76]*tmp[198]+tmp[77]*tmp[197]+tmp[78]*tmp[196]+tmp[79]*tmp[195]+tmp[80]*tmp[194]+tmp[81]*tmp[193]+tmp[82]*tmp[192]+tmp[83]*tmp[191]+tmp[84]*tmp[190]+tmp[85]*tmp[189]+tmp[86]*tmp[188]+tmp[87]*tmp[187]+tmp[88]*tmp[186]+tmp[89]*tmp[185]+tmp[90]*tmp[184]+tmp[91]*tmp[183]+tmp[92]*tmp[182]+tmp[93]*tmp[181]+tmp[94]*tmp[180]+tmp[95]*tmp[179]+tmp[96]*tmp[178]+tmp[97]*tmp[177]+tmp[98]*tmp[176]+tmp[99]*tmp[175];
				ans[175]<=tmp[76]*tmp[199]+tmp[77]*tmp[198]+tmp[78]*tmp[197]+tmp[79]*tmp[196]+tmp[80]*tmp[195]+tmp[81]*tmp[194]+tmp[82]*tmp[193]+tmp[83]*tmp[192]+tmp[84]*tmp[191]+tmp[85]*tmp[190]+tmp[86]*tmp[189]+tmp[87]*tmp[188]+tmp[88]*tmp[187]+tmp[89]*tmp[186]+tmp[90]*tmp[185]+tmp[91]*tmp[184]+tmp[92]*tmp[183]+tmp[93]*tmp[182]+tmp[94]*tmp[181]+tmp[95]*tmp[180]+tmp[96]*tmp[179]+tmp[97]*tmp[178]+tmp[98]*tmp[177]+tmp[99]*tmp[176];
				ans[176]<=tmp[77]*tmp[199]+tmp[78]*tmp[198]+tmp[79]*tmp[197]+tmp[80]*tmp[196]+tmp[81]*tmp[195]+tmp[82]*tmp[194]+tmp[83]*tmp[193]+tmp[84]*tmp[192]+tmp[85]*tmp[191]+tmp[86]*tmp[190]+tmp[87]*tmp[189]+tmp[88]*tmp[188]+tmp[89]*tmp[187]+tmp[90]*tmp[186]+tmp[91]*tmp[185]+tmp[92]*tmp[184]+tmp[93]*tmp[183]+tmp[94]*tmp[182]+tmp[95]*tmp[181]+tmp[96]*tmp[180]+tmp[97]*tmp[179]+tmp[98]*tmp[178]+tmp[99]*tmp[177];
				ans[177]<=tmp[78]*tmp[199]+tmp[79]*tmp[198]+tmp[80]*tmp[197]+tmp[81]*tmp[196]+tmp[82]*tmp[195]+tmp[83]*tmp[194]+tmp[84]*tmp[193]+tmp[85]*tmp[192]+tmp[86]*tmp[191]+tmp[87]*tmp[190]+tmp[88]*tmp[189]+tmp[89]*tmp[188]+tmp[90]*tmp[187]+tmp[91]*tmp[186]+tmp[92]*tmp[185]+tmp[93]*tmp[184]+tmp[94]*tmp[183]+tmp[95]*tmp[182]+tmp[96]*tmp[181]+tmp[97]*tmp[180]+tmp[98]*tmp[179]+tmp[99]*tmp[178];
				ans[178]<=tmp[79]*tmp[199]+tmp[80]*tmp[198]+tmp[81]*tmp[197]+tmp[82]*tmp[196]+tmp[83]*tmp[195]+tmp[84]*tmp[194]+tmp[85]*tmp[193]+tmp[86]*tmp[192]+tmp[87]*tmp[191]+tmp[88]*tmp[190]+tmp[89]*tmp[189]+tmp[90]*tmp[188]+tmp[91]*tmp[187]+tmp[92]*tmp[186]+tmp[93]*tmp[185]+tmp[94]*tmp[184]+tmp[95]*tmp[183]+tmp[96]*tmp[182]+tmp[97]*tmp[181]+tmp[98]*tmp[180]+tmp[99]*tmp[179];
				ans[179]<=tmp[80]*tmp[199]+tmp[81]*tmp[198]+tmp[82]*tmp[197]+tmp[83]*tmp[196]+tmp[84]*tmp[195]+tmp[85]*tmp[194]+tmp[86]*tmp[193]+tmp[87]*tmp[192]+tmp[88]*tmp[191]+tmp[89]*tmp[190]+tmp[90]*tmp[189]+tmp[91]*tmp[188]+tmp[92]*tmp[187]+tmp[93]*tmp[186]+tmp[94]*tmp[185]+tmp[95]*tmp[184]+tmp[96]*tmp[183]+tmp[97]*tmp[182]+tmp[98]*tmp[181]+tmp[99]*tmp[180];
				ans[180]<=tmp[81]*tmp[199]+tmp[82]*tmp[198]+tmp[83]*tmp[197]+tmp[84]*tmp[196]+tmp[85]*tmp[195]+tmp[86]*tmp[194]+tmp[87]*tmp[193]+tmp[88]*tmp[192]+tmp[89]*tmp[191]+tmp[90]*tmp[190]+tmp[91]*tmp[189]+tmp[92]*tmp[188]+tmp[93]*tmp[187]+tmp[94]*tmp[186]+tmp[95]*tmp[185]+tmp[96]*tmp[184]+tmp[97]*tmp[183]+tmp[98]*tmp[182]+tmp[99]*tmp[181];
				ans[181]<=tmp[82]*tmp[199]+tmp[83]*tmp[198]+tmp[84]*tmp[197]+tmp[85]*tmp[196]+tmp[86]*tmp[195]+tmp[87]*tmp[194]+tmp[88]*tmp[193]+tmp[89]*tmp[192]+tmp[90]*tmp[191]+tmp[91]*tmp[190]+tmp[92]*tmp[189]+tmp[93]*tmp[188]+tmp[94]*tmp[187]+tmp[95]*tmp[186]+tmp[96]*tmp[185]+tmp[97]*tmp[184]+tmp[98]*tmp[183]+tmp[99]*tmp[182];
				ans[182]<=tmp[83]*tmp[199]+tmp[84]*tmp[198]+tmp[85]*tmp[197]+tmp[86]*tmp[196]+tmp[87]*tmp[195]+tmp[88]*tmp[194]+tmp[89]*tmp[193]+tmp[90]*tmp[192]+tmp[91]*tmp[191]+tmp[92]*tmp[190]+tmp[93]*tmp[189]+tmp[94]*tmp[188]+tmp[95]*tmp[187]+tmp[96]*tmp[186]+tmp[97]*tmp[185]+tmp[98]*tmp[184]+tmp[99]*tmp[183];
				ans[183]<=tmp[84]*tmp[199]+tmp[85]*tmp[198]+tmp[86]*tmp[197]+tmp[87]*tmp[196]+tmp[88]*tmp[195]+tmp[89]*tmp[194]+tmp[90]*tmp[193]+tmp[91]*tmp[192]+tmp[92]*tmp[191]+tmp[93]*tmp[190]+tmp[94]*tmp[189]+tmp[95]*tmp[188]+tmp[96]*tmp[187]+tmp[97]*tmp[186]+tmp[98]*tmp[185]+tmp[99]*tmp[184];
				ans[184]<=tmp[85]*tmp[199]+tmp[86]*tmp[198]+tmp[87]*tmp[197]+tmp[88]*tmp[196]+tmp[89]*tmp[195]+tmp[90]*tmp[194]+tmp[91]*tmp[193]+tmp[92]*tmp[192]+tmp[93]*tmp[191]+tmp[94]*tmp[190]+tmp[95]*tmp[189]+tmp[96]*tmp[188]+tmp[97]*tmp[187]+tmp[98]*tmp[186]+tmp[99]*tmp[185];
				ans[185]<=tmp[86]*tmp[199]+tmp[87]*tmp[198]+tmp[88]*tmp[197]+tmp[89]*tmp[196]+tmp[90]*tmp[195]+tmp[91]*tmp[194]+tmp[92]*tmp[193]+tmp[93]*tmp[192]+tmp[94]*tmp[191]+tmp[95]*tmp[190]+tmp[96]*tmp[189]+tmp[97]*tmp[188]+tmp[98]*tmp[187]+tmp[99]*tmp[186];
				ans[186]<=tmp[87]*tmp[199]+tmp[88]*tmp[198]+tmp[89]*tmp[197]+tmp[90]*tmp[196]+tmp[91]*tmp[195]+tmp[92]*tmp[194]+tmp[93]*tmp[193]+tmp[94]*tmp[192]+tmp[95]*tmp[191]+tmp[96]*tmp[190]+tmp[97]*tmp[189]+tmp[98]*tmp[188]+tmp[99]*tmp[187];
				ans[187]<=tmp[88]*tmp[199]+tmp[89]*tmp[198]+tmp[90]*tmp[197]+tmp[91]*tmp[196]+tmp[92]*tmp[195]+tmp[93]*tmp[194]+tmp[94]*tmp[193]+tmp[95]*tmp[192]+tmp[96]*tmp[191]+tmp[97]*tmp[190]+tmp[98]*tmp[189]+tmp[99]*tmp[188];
				ans[188]<=tmp[89]*tmp[199]+tmp[90]*tmp[198]+tmp[91]*tmp[197]+tmp[92]*tmp[196]+tmp[93]*tmp[195]+tmp[94]*tmp[194]+tmp[95]*tmp[193]+tmp[96]*tmp[192]+tmp[97]*tmp[191]+tmp[98]*tmp[190]+tmp[99]*tmp[189];
				ans[189]<=tmp[90]*tmp[199]+tmp[91]*tmp[198]+tmp[92]*tmp[197]+tmp[93]*tmp[196]+tmp[94]*tmp[195]+tmp[95]*tmp[194]+tmp[96]*tmp[193]+tmp[97]*tmp[192]+tmp[98]*tmp[191]+tmp[99]*tmp[190];
				ans[190]<=tmp[91]*tmp[199]+tmp[92]*tmp[198]+tmp[93]*tmp[197]+tmp[94]*tmp[196]+tmp[95]*tmp[195]+tmp[96]*tmp[194]+tmp[97]*tmp[193]+tmp[98]*tmp[192]+tmp[99]*tmp[191];
				ans[191]<=tmp[92]*tmp[199]+tmp[93]*tmp[198]+tmp[94]*tmp[197]+tmp[95]*tmp[196]+tmp[96]*tmp[195]+tmp[97]*tmp[194]+tmp[98]*tmp[193]+tmp[99]*tmp[192];
				ans[192]<=tmp[93]*tmp[199]+tmp[94]*tmp[198]+tmp[95]*tmp[197]+tmp[96]*tmp[196]+tmp[97]*tmp[195]+tmp[98]*tmp[194]+tmp[99]*tmp[193];
				ans[193]<=tmp[94]*tmp[199]+tmp[95]*tmp[198]+tmp[96]*tmp[197]+tmp[97]*tmp[196]+tmp[98]*tmp[195]+tmp[99]*tmp[194];
				ans[194]<=tmp[95]*tmp[199]+tmp[96]*tmp[198]+tmp[97]*tmp[197]+tmp[98]*tmp[196]+tmp[99]*tmp[195];
				ans[195]<=tmp[96]*tmp[199]+tmp[97]*tmp[198]+tmp[98]*tmp[197]+tmp[99]*tmp[196];
				ans[196]<=tmp[97]*tmp[199]+tmp[98]*tmp[198]+tmp[99]*tmp[197];
				ans[197]<=tmp[98]*tmp[199]+tmp[99]*tmp[198];
				ans[198]<=tmp[99]*tmp[199];
                state<=READY_WRITE;
            end
            else if (state == READY_WRITE)
            begin
                r_write_addr<=write_base;
                r_write_size<=read_size_input;
                r_write_data <= ans[write_cnt[7:0]];
                r_write_enable<=1;
                state<=WAIT_WRITE;
            end
            else if (state == WAIT_WRITE)
            begin
                r_finish_write<=0;
                if (write_ready == 1)
                begin
                    state<=DEAL_WRITE;
                end
            end
            else if (state == DEAL_WRITE)
            begin
                if (write_cnt + 1 < num_read)
                begin
                    r_finish_write<=1;
                    write_cnt<=write_cnt+1;
                    r_write_data<=ans[write_cnt[7:0]];
                    r_write_addr<=r_write_addr+write_size;
                    state<=WAIT_WRITE;
                end
                else
                begin
                    r_finish_write<=0;
                    r_write_enable<=0;
                    state<=SUSPEND;
                    r_done<=1;
                end
            end
			
        end
    end
endmodule
